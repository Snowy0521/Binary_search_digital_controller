// Created by ihdl
module FIR_Filter ( CLK_Filter, input_data, rst_n, output_data );
  input [7:0] input_data;
  output [19:0] output_data;
  input CLK_Filter, rst_n;
  wire   N1, N2, N3, N4, N5, N6, N7, N8, N10, N11, N12, N13, N14, N15, N16,
         N17, N19, N20, N21, N22, N23, N24, N25, N26, N28, N29, N30, N31, N32,
         N33, N34, N35, N37, N38, N39, N40, N41, N42, N43, N44, N46, N47, N48,
         N49, N50, N51, N52, N53, N55, N56, N57, N58, N59, N60, N61, N62, N64,
         N65, N66, N67, N68, N69, N70, N71, N73, N74, N75, N76, N77, N78, N79,
         N80, N82, N83, N84, N85, N86, N87, N88, N89, N91, N92, N93, N94, N95,
         N96, N97, N98, N101, N102, N103, N104, N105, N106, N107, N108, N109,
         N110, N111, N112, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N144, N145, N146,
         N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N158,
         N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N398, N399, N400, N401, N402,
         N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413,
         N414, N415, intadd_0_A_17_, intadd_0_A_16_, intadd_0_A_15_,
         intadd_0_A_14_, intadd_0_A_13_, intadd_0_A_12_, intadd_0_A_11_,
         intadd_0_A_10_, intadd_0_A_9_, intadd_0_A_8_, intadd_0_A_7_,
         intadd_0_A_6_, intadd_0_A_5_, intadd_0_A_4_, intadd_0_A_3_,
         intadd_0_A_2_, intadd_0_A_1_, intadd_0_B_5_, intadd_0_B_3_,
         intadd_0_B_2_, intadd_0_B_1_, intadd_0_n18, intadd_0_n17,
         intadd_0_n16, intadd_0_n15, intadd_0_n14, intadd_0_n13, intadd_0_n12,
         intadd_0_n11, intadd_0_n10, intadd_0_n9, intadd_0_n8, intadd_0_n7,
         intadd_0_n6, intadd_0_n5, intadd_0_n4, intadd_0_n3, intadd_0_n2,
         intadd_0_n1, intadd_1_A_8_, intadd_1_A_7_, intadd_1_A_6_,
         intadd_1_A_5_, intadd_1_A_4_, intadd_1_A_3_, intadd_1_A_2_,
         intadd_1_A_1_, intadd_1_B_9_, intadd_1_B_8_, intadd_1_B_7_,
         intadd_1_B_6_, intadd_1_B_5_, intadd_1_B_4_, intadd_1_B_3_,
         intadd_1_B_2_, intadd_1_B_1_, intadd_1_B_0_, intadd_1_CI,
         intadd_1_n10, intadd_1_n9, intadd_1_n8, intadd_1_n7, intadd_1_n6,
         intadd_1_n5, intadd_1_n4, intadd_1_n3, intadd_1_n2, intadd_1_n1,
         intadd_2_A_7_, intadd_2_A_6_, intadd_2_A_5_, intadd_2_A_4_,
         intadd_2_A_3_, intadd_2_B_7_, intadd_2_B_6_, intadd_2_B_5_,
         intadd_2_B_4_, intadd_2_B_3_, intadd_2_B_2_, intadd_2_B_1_,
         intadd_2_B_0_, intadd_2_CI, intadd_2_SUM_7_, intadd_2_SUM_6_,
         intadd_2_SUM_5_, intadd_2_SUM_4_, intadd_2_SUM_3_, intadd_2_SUM_2_,
         intadd_2_SUM_1_, intadd_2_SUM_0_, intadd_2_n8, intadd_2_n7,
         intadd_2_n6, intadd_2_n5, intadd_2_n4, intadd_2_n3, intadd_2_n2,
         intadd_2_n1, intadd_3_A_6_, intadd_3_A_5_, intadd_3_A_4_,
         intadd_3_A_3_, intadd_3_A_2_, intadd_3_A_1_, intadd_3_B_6_,
         intadd_3_B_5_, intadd_3_B_4_, intadd_3_B_3_, intadd_3_B_2_,
         intadd_3_B_1_, intadd_3_B_0_, intadd_3_CI, intadd_3_SUM_6_,
         intadd_3_SUM_5_, intadd_3_SUM_4_, intadd_3_SUM_3_, intadd_3_SUM_2_,
         intadd_3_SUM_1_, intadd_3_SUM_0_, intadd_3_n7, intadd_3_n6,
         intadd_3_n5, intadd_3_n4, intadd_3_n3, intadd_3_n2, intadd_3_n1,
         intadd_4_A_6_, intadd_4_A_5_, intadd_4_A_4_, intadd_4_A_3_,
         intadd_4_A_2_, intadd_4_A_1_, intadd_4_B_6_, intadd_4_B_5_,
         intadd_4_B_4_, intadd_4_B_3_, intadd_4_B_2_, intadd_4_B_1_,
         intadd_4_B_0_, intadd_4_CI, intadd_4_n7, intadd_4_n6, intadd_4_n5,
         intadd_4_n4, intadd_4_n3, intadd_4_n2, intadd_4_n1, intadd_5_CI,
         intadd_5_n7, intadd_5_n6, intadd_5_n5, intadd_5_n4, intadd_5_n3,
         intadd_5_n2, intadd_5_n1, intadd_6_CI, intadd_6_n7, intadd_6_n6,
         intadd_6_n5, intadd_6_n4, intadd_6_n3, intadd_6_n2, intadd_6_n1,
         intadd_7_CI, intadd_7_n7, intadd_7_n6, intadd_7_n5, intadd_7_n4,
         intadd_7_n3, intadd_7_n2, intadd_7_n1, intadd_8_CI, intadd_8_n7,
         intadd_8_n6, intadd_8_n5, intadd_8_n4, intadd_8_n3, intadd_8_n2,
         intadd_8_n1, intadd_9_CI, intadd_9_n7, intadd_9_n6, intadd_9_n5,
         intadd_9_n4, intadd_9_n3, intadd_9_n2, intadd_9_n1, intadd_10_CI,
         intadd_10_n7, intadd_10_n6, intadd_10_n5, intadd_10_n4, intadd_10_n3,
         intadd_10_n2, intadd_10_n1, intadd_11_CI, intadd_11_n7, intadd_11_n6,
         intadd_11_n5, intadd_11_n4, intadd_11_n3, intadd_11_n2, intadd_11_n1,
         intadd_12_CI, intadd_12_n7, intadd_12_n6, intadd_12_n5, intadd_12_n4,
         intadd_12_n3, intadd_12_n2, intadd_12_n1, intadd_13_CI, intadd_13_n7,
         intadd_13_n6, intadd_13_n5, intadd_13_n4, intadd_13_n3, intadd_13_n2,
         intadd_13_n1, intadd_14_CI, intadd_14_n7, intadd_14_n6, intadd_14_n5,
         intadd_14_n4, intadd_14_n3, intadd_14_n2, intadd_14_n1, intadd_15_CI,
         intadd_15_n7, intadd_15_n6, intadd_15_n5, intadd_15_n4, intadd_15_n3,
         intadd_15_n2, intadd_15_n1, intadd_16_CI, intadd_16_n6, intadd_16_n5,
         intadd_16_n4, intadd_16_n3, intadd_16_n2, intadd_16_n1,
         intadd_17_A_4_, intadd_17_A_3_, intadd_17_A_2_, intadd_17_A_1_,
         intadd_17_B_3_, intadd_17_B_2_, intadd_17_B_1_, intadd_17_SUM_3_,
         intadd_17_SUM_2_, intadd_17_SUM_1_, intadd_17_SUM_0_, intadd_17_n5,
         intadd_17_n4, intadd_17_n3, intadd_17_n2, intadd_17_n1,
         intadd_18_A_4_, intadd_18_A_3_, intadd_18_A_1_, intadd_18_B_3_,
         intadd_18_B_2_, intadd_18_B_1_, intadd_18_SUM_3_, intadd_18_SUM_2_,
         intadd_18_SUM_1_, intadd_18_SUM_0_, intadd_18_n5, intadd_18_n4,
         intadd_18_n3, intadd_18_n2, intadd_18_n1, intadd_19_A_3_,
         intadd_19_A_2_, intadd_19_A_1_, intadd_19_B_2_, intadd_19_B_1_,
         intadd_19_SUM_3_, intadd_19_SUM_2_, intadd_19_SUM_1_,
         intadd_19_SUM_0_, intadd_19_n5, intadd_19_n4, intadd_19_n3,
         intadd_19_n2, intadd_19_n1, intadd_20_A_3_, intadd_20_A_2_,
         intadd_20_A_1_, intadd_20_B_2_, intadd_20_B_1_, intadd_20_SUM_3_,
         intadd_20_SUM_2_, intadd_20_SUM_1_, intadd_20_SUM_0_, intadd_20_n5,
         intadd_20_n4, intadd_20_n3, intadd_20_n2, intadd_20_n1,
         intadd_21_A_3_, intadd_21_A_2_, intadd_21_A_1_, intadd_21_B_2_,
         intadd_21_B_1_, intadd_21_SUM_3_, intadd_21_SUM_2_, intadd_21_SUM_1_,
         intadd_21_SUM_0_, intadd_21_n5, intadd_21_n4, intadd_21_n3,
         intadd_21_n2, intadd_21_n1, intadd_22_A_3_, intadd_22_B_2_,
         intadd_22_B_1_, intadd_22_SUM_3_, intadd_22_SUM_2_, intadd_22_SUM_1_,
         intadd_22_SUM_0_, intadd_22_n5, intadd_22_n4, intadd_22_n3,
         intadd_22_n2, intadd_22_n1, intadd_23_A_3_, intadd_23_B_2_,
         intadd_23_SUM_3_, intadd_23_SUM_2_, intadd_23_SUM_1_,
         intadd_23_SUM_0_, intadd_23_n5, intadd_23_n4, intadd_23_n3,
         intadd_23_n2, intadd_23_n1, intadd_24_A_3_, intadd_24_A_2_,
         intadd_24_B_1_, intadd_24_SUM_3_, intadd_24_SUM_2_, intadd_24_SUM_1_,
         intadd_24_SUM_0_, intadd_24_n5, intadd_24_n4, intadd_24_n3,
         intadd_24_n2, intadd_24_n1, intadd_25_A_1_, intadd_25_A_0_,
         intadd_25_B_4_, intadd_25_B_3_, intadd_25_B_2_, intadd_25_CI,
         intadd_25_SUM_4_, intadd_25_SUM_3_, intadd_25_SUM_2_,
         intadd_25_SUM_1_, intadd_25_SUM_0_, intadd_25_n5, intadd_25_n4,
         intadd_25_n3, intadd_25_n2, intadd_25_n1, intadd_26_A_3_,
         intadd_26_A_2_, intadd_26_A_1_, intadd_26_B_3_, intadd_26_B_2_,
         intadd_26_B_1_, intadd_26_SUM_2_, intadd_26_SUM_1_, intadd_26_SUM_0_,
         intadd_26_n4, intadd_26_n3, intadd_26_n2, intadd_26_n1,
         intadd_27_A_2_, intadd_27_A_1_, intadd_27_B_3_, intadd_27_B_2_,
         intadd_27_B_1_, intadd_27_SUM_2_, intadd_27_SUM_1_, intadd_27_SUM_0_,
         intadd_27_n4, intadd_27_n3, intadd_27_n2, intadd_27_n1,
         intadd_28_A_2_, intadd_28_A_1_, intadd_28_B_1_, intadd_28_SUM_2_,
         intadd_28_SUM_1_, intadd_28_SUM_0_, intadd_28_n4, intadd_28_n3,
         intadd_28_n2, intadd_28_n1, intadd_29_A_1_, intadd_29_B_1_,
         intadd_29_SUM_2_, intadd_29_SUM_1_, intadd_29_SUM_0_, intadd_29_n4,
         intadd_29_n3, intadd_29_n2, intadd_29_n1, intadd_30_B_3_,
         intadd_30_B_2_, intadd_30_B_1_, intadd_30_B_0_, intadd_30_CI,
         intadd_30_SUM_3_, intadd_30_SUM_2_, intadd_30_SUM_1_,
         intadd_30_SUM_0_, intadd_30_n4, intadd_30_n3, intadd_30_n2,
         intadd_30_n1, intadd_31_A_3_, intadd_31_A_2_, intadd_31_A_1_,
         intadd_31_B_3_, intadd_31_B_2_, intadd_31_B_1_, intadd_31_CI,
         intadd_31_SUM_0_, intadd_31_n4, intadd_31_n3, intadd_31_n2,
         intadd_31_n1, intadd_32_A_3_, intadd_32_A_2_, intadd_32_A_1_,
         intadd_32_B_3_, intadd_32_B_2_, intadd_32_B_1_, intadd_32_B_0_,
         intadd_32_CI, intadd_32_SUM_3_, intadd_32_SUM_2_, intadd_32_SUM_1_,
         intadd_32_SUM_0_, intadd_32_n4, intadd_32_n3, intadd_32_n2,
         intadd_32_n1, intadd_33_A_2_, intadd_33_SUM_0_, intadd_33_n3,
         intadd_33_n2, intadd_33_n1, intadd_34_A_1_, intadd_34_B_2_,
         intadd_34_B_1_, intadd_34_SUM_0_, intadd_34_n3, intadd_34_n2,
         intadd_34_n1, intadd_35_A_1_, intadd_35_B_2_, intadd_35_B_1_,
         intadd_35_n3, intadd_35_n2, intadd_35_n1, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158;
  wire   [175:0] shift_regs;
  wire   [140:0] order;
  wire   [88:0] add_regs;

  DFQRM1SA output_data_reg_4_ ( .D(N402), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[4]) );
  DFQRM1SA order_reg_9__5_ ( .D(N210), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[121]) );
  DFQRM1SA order_reg_8__5_ ( .D(N194), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[106]) );
  DFQRM1SA order_reg_7__6_ ( .D(N179), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[91]) );
  DFQRM1SA order_reg_6__7_ ( .D(N164), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[76]) );
  DFQRM1SA order_reg_5__6_ ( .D(N148), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[61]) );
  DFQRM1SA order_reg_4__4_ ( .D(N131), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[46]) );
  DFQRM1SA order_reg_3__3_ ( .D(N116), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[31]) );
  DFQRM1SA order_reg_10__15_ ( .D(add_regs[88]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[140]) );
  DFQRM1SA add_regs_reg_10__0_ ( .D(N91), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[80]) );
  DFQRM1SA add_regs_reg_8__4_ ( .D(N77), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[68]) );
  DFQRM1SA add_regs_reg_6__7_ ( .D(N62), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[55]) );
  DFQRM1SA add_regs_reg_5__1_ ( .D(N47), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[41]) );
  DFQRM1SA add_regs_reg_3__4_ ( .D(N32), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[28]) );
  DFQRM1SA add_regs_reg_2__3_ ( .D(N22), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[19]) );
  DFQRM1SA add_regs_reg_1__1_ ( .D(N11), .CK(CLK_Filter), .RB(rst_n), .Q(N102)
         );
  DFQRM1SA order_reg_0__3_ ( .D(add_regs[2]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[2]) );
  DFQRM1SA shift_regs_reg_10__7_ ( .D(shift_regs[79]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[87]) );
  DFQRM1SA shift_regs_reg_3__6_ ( .D(shift_regs[22]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[30]) );
  DFQRM1SA shift_regs_reg_18__6_ ( .D(shift_regs[142]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[150]) );
  DFQRM1SA shift_regs_reg_11__5_ ( .D(shift_regs[85]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[93]) );
  DFQRM1SA shift_regs_reg_4__4_ ( .D(shift_regs[28]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[36]) );
  DFQRM1SA shift_regs_reg_19__4_ ( .D(shift_regs[148]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[156]) );
  DFQRM1SA shift_regs_reg_12__3_ ( .D(shift_regs[91]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[99]) );
  DFQRM1SA shift_regs_reg_5__2_ ( .D(shift_regs[34]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[42]) );
  DFQRM1SA shift_regs_reg_20__2_ ( .D(shift_regs[154]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[162]) );
  DFQRM1SA shift_regs_reg_13__1_ ( .D(shift_regs[97]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[105]) );
  DFQRM1SA shift_regs_reg_6__0_ ( .D(shift_regs[40]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[48]) );
  DFQRM1SA shift_regs_reg_21__0_ ( .D(shift_regs[160]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[168]) );
  DFQRM1SA output_data_reg_18_ ( .D(intadd_0_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(output_data[18]) );
  DFQRM1SA output_data_reg_17_ ( .D(N415), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[17]) );
  DFQRM1SA output_data_reg_16_ ( .D(N414), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[16]) );
  DFQRM1SA output_data_reg_15_ ( .D(N413), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[15]) );
  DFQRM1SA output_data_reg_14_ ( .D(N412), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[14]) );
  DFQRM1SA output_data_reg_13_ ( .D(N411), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[13]) );
  DFQRM1SA output_data_reg_12_ ( .D(N410), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[12]) );
  DFQRM1SA output_data_reg_11_ ( .D(N409), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[11]) );
  DFQRM1SA output_data_reg_10_ ( .D(N408), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[10]) );
  DFQRM1SA output_data_reg_9_ ( .D(N407), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[9]) );
  DFQRM1SA output_data_reg_8_ ( .D(N406), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[8]) );
  DFQRM1SA output_data_reg_7_ ( .D(N405), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[7]) );
  DFQRM1SA output_data_reg_6_ ( .D(N404), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[6]) );
  DFQRM1SA output_data_reg_5_ ( .D(N403), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[5]) );
  DFQRM1SA output_data_reg_3_ ( .D(N401), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[3]) );
  DFQRM1SA output_data_reg_2_ ( .D(N400), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[2]) );
  DFQRM1SA output_data_reg_1_ ( .D(N399), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[1]) );
  DFQRM1SA output_data_reg_0_ ( .D(N398), .CK(CLK_Filter), .RB(rst_n), .Q(
        output_data[0]) );
  DFQRM1SA order_reg_9__15_ ( .D(N220), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[131]) );
  DFQRM1SA order_reg_9__14_ ( .D(N219), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[130]) );
  DFQRM1SA order_reg_9__13_ ( .D(N218), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[129]) );
  DFQRM1SA order_reg_9__12_ ( .D(N217), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[128]) );
  DFQRM1SA order_reg_9__11_ ( .D(N216), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[127]) );
  DFQRM1SA order_reg_9__10_ ( .D(N215), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[126]) );
  DFQRM1SA order_reg_9__9_ ( .D(N214), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[125]) );
  DFQRM1SA order_reg_9__8_ ( .D(N213), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[124]) );
  DFQRM1SA order_reg_9__7_ ( .D(N212), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[123]) );
  DFQRM1SA order_reg_9__6_ ( .D(N211), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[122]) );
  DFQRM1SA order_reg_9__4_ ( .D(N209), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[120]) );
  DFQRM1SA order_reg_9__3_ ( .D(N208), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[119]) );
  DFQRM1SA order_reg_8__15_ ( .D(N204), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[116]) );
  DFQRM1SA order_reg_8__14_ ( .D(N203), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[115]) );
  DFQRM1SA order_reg_8__13_ ( .D(N202), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[114]) );
  DFQRM1SA order_reg_8__12_ ( .D(N201), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[113]) );
  DFQRM1SA order_reg_8__11_ ( .D(N200), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[112]) );
  DFQRM1SA order_reg_8__10_ ( .D(N199), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[111]) );
  DFQRM1SA order_reg_8__9_ ( .D(N198), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[110]) );
  DFQRM1SA order_reg_8__8_ ( .D(N197), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[109]) );
  DFQRM1SA order_reg_8__7_ ( .D(N196), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[108]) );
  DFQRM1SA order_reg_8__6_ ( .D(N195), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[107]) );
  DFQRM1SA order_reg_8__4_ ( .D(N193), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[105]) );
  DFQRM1SA order_reg_8__3_ ( .D(N192), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[104]) );
  DFQRM1SA order_reg_8__2_ ( .D(N191), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[103]) );
  DFQRM1SA order_reg_8__1_ ( .D(N190), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[102]) );
  DFQRM1SA order_reg_7__15_ ( .D(N188), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[100]) );
  DFQRM1SA order_reg_7__14_ ( .D(N187), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[99]) );
  DFQRM1SA order_reg_7__13_ ( .D(N186), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[98]) );
  DFQRM1SA order_reg_7__12_ ( .D(N185), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[97]) );
  DFQRM1SA order_reg_7__11_ ( .D(N184), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[96]) );
  DFQRM1SA order_reg_7__10_ ( .D(N183), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[95]) );
  DFQRM1SA order_reg_7__9_ ( .D(N182), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[94]) );
  DFQRM1SA order_reg_7__8_ ( .D(N181), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[93]) );
  DFQRM1SA order_reg_7__7_ ( .D(N180), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[92]) );
  DFQRM1SA order_reg_7__5_ ( .D(N178), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[90]) );
  DFQRM1SA order_reg_7__4_ ( .D(N177), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[89]) );
  DFQRM1SA order_reg_7__3_ ( .D(N176), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[88]) );
  DFQRM1SA order_reg_7__2_ ( .D(N175), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[87]) );
  DFQRM1SA order_reg_7__1_ ( .D(N174), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[86]) );
  DFQRM1SA order_reg_6__15_ ( .D(N172), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[84]) );
  DFQRM1SA order_reg_6__14_ ( .D(N171), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[83]) );
  DFQRM1SA order_reg_6__13_ ( .D(N170), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[82]) );
  DFQRM1SA order_reg_6__12_ ( .D(N169), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[81]) );
  DFQRM1SA order_reg_6__11_ ( .D(N168), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[80]) );
  DFQRM1SA order_reg_6__10_ ( .D(N167), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[79]) );
  DFQRM1SA order_reg_6__9_ ( .D(N166), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[78]) );
  DFQRM1SA order_reg_6__8_ ( .D(N165), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[77]) );
  DFQRM1SA order_reg_6__6_ ( .D(N163), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[75]) );
  DFQRM1SA order_reg_6__5_ ( .D(N162), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[74]) );
  DFQRM1SA order_reg_6__4_ ( .D(N161), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[73]) );
  DFQRM1SA order_reg_6__3_ ( .D(N160), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[72]) );
  DFQRM1SA order_reg_6__2_ ( .D(N159), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[71]) );
  DFQRM1SA order_reg_5__14_ ( .D(N156), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[69]) );
  DFQRM1SA order_reg_5__13_ ( .D(N155), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[68]) );
  DFQRM1SA order_reg_5__12_ ( .D(N154), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[67]) );
  DFQRM1SA order_reg_5__11_ ( .D(N153), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[66]) );
  DFQRM1SA order_reg_5__10_ ( .D(N152), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[65]) );
  DFQRM1SA order_reg_5__9_ ( .D(N151), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[64]) );
  DFQRM1SA order_reg_5__8_ ( .D(N150), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[63]) );
  DFQRM1SA order_reg_5__7_ ( .D(N149), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[62]) );
  DFQRM1SA order_reg_5__5_ ( .D(N147), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[60]) );
  DFQRM1SA order_reg_5__4_ ( .D(N146), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[59]) );
  DFQRM1SA order_reg_5__3_ ( .D(N145), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[58]) );
  DFQRM1SA order_reg_4__14_ ( .D(N141), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[56]) );
  DFQRM1SA order_reg_4__13_ ( .D(N140), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[55]) );
  DFQRM1SA order_reg_4__12_ ( .D(N139), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[54]) );
  DFQRM1SA order_reg_4__11_ ( .D(N138), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[53]) );
  DFQRM1SA order_reg_4__10_ ( .D(N137), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[52]) );
  DFQRM1SA order_reg_4__9_ ( .D(N136), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[51]) );
  DFQRM1SA order_reg_4__8_ ( .D(N135), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[50]) );
  DFQRM1SA order_reg_4__7_ ( .D(N134), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[49]) );
  DFQRM1SA order_reg_4__6_ ( .D(N133), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[48]) );
  DFQRM1SA order_reg_4__5_ ( .D(N132), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[47]) );
  DFQRM1SA order_reg_4__3_ ( .D(N130), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[45]) );
  DFQRM1SA order_reg_4__2_ ( .D(N129), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[44]) );
  DFQRM1SA order_reg_4__1_ ( .D(N128), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[43]) );
  DFQRM1SA order_reg_3__13_ ( .D(N126), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[41]) );
  DFQRM1SA order_reg_3__12_ ( .D(N125), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[40]) );
  DFQRM1SA order_reg_3__11_ ( .D(N124), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[39]) );
  DFQRM1SA order_reg_3__10_ ( .D(N123), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[38]) );
  DFQRM1SA order_reg_3__9_ ( .D(N122), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[37]) );
  DFQRM1SA order_reg_3__8_ ( .D(N121), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[36]) );
  DFQRM1SA order_reg_3__7_ ( .D(N120), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[35]) );
  DFQRM1SA order_reg_3__6_ ( .D(N119), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[34]) );
  DFQRM1SA order_reg_3__5_ ( .D(N118), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[33]) );
  DFQRM1SA order_reg_3__4_ ( .D(N117), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[32]) );
  DFQRM1SA order_reg_1__12_ ( .D(N112), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[20]) );
  DFQRM1SA order_reg_1__11_ ( .D(N111), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[19]) );
  DFQRM1SA order_reg_1__10_ ( .D(N110), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[18]) );
  DFQRM1SA order_reg_1__9_ ( .D(N109), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[17]) );
  DFQRM1SA order_reg_1__8_ ( .D(N108), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[16]) );
  DFQRM1SA order_reg_1__7_ ( .D(N107), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[15]) );
  DFQRM1SA order_reg_1__6_ ( .D(N106), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[14]) );
  DFQRM1SA order_reg_1__5_ ( .D(N105), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[13]) );
  DFQRM1SA order_reg_1__4_ ( .D(N104), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[12]) );
  DFQRM1SA order_reg_1__3_ ( .D(N103), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[11]) );
  DFQRM1SA add_regs_reg_10__8_ ( .D(intadd_5_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[88]) );
  DFQRM1SA add_regs_reg_10__7_ ( .D(N98), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[87]) );
  DFQRM1SA add_regs_reg_10__6_ ( .D(N97), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[86]) );
  DFQRM1SA add_regs_reg_10__5_ ( .D(N96), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[85]) );
  DFQRM1SA add_regs_reg_10__4_ ( .D(N95), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[84]) );
  DFQRM1SA add_regs_reg_10__3_ ( .D(N94), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[83]) );
  DFQRM1SA add_regs_reg_10__2_ ( .D(N93), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[82]) );
  DFQRM1SA add_regs_reg_10__1_ ( .D(N92), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[81]) );
  DFQRM1SA add_regs_reg_9__8_ ( .D(intadd_6_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[79]) );
  DFQRM1SA add_regs_reg_9__7_ ( .D(N89), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[78]) );
  DFQRM1SA add_regs_reg_9__6_ ( .D(N88), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[77]) );
  DFQRM1SA add_regs_reg_9__5_ ( .D(N87), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[76]) );
  DFQRM1SA add_regs_reg_9__4_ ( .D(N86), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[75]) );
  DFQRM1SA add_regs_reg_9__3_ ( .D(N85), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[74]) );
  DFQRM1SA add_regs_reg_9__2_ ( .D(N84), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[73]) );
  DFQRM1SA add_regs_reg_9__1_ ( .D(N83), .CK(CLK_Filter), .RB(rst_n), .Q(N207)
         );
  DFQRM1SA add_regs_reg_9__0_ ( .D(N82), .CK(CLK_Filter), .RB(rst_n), .Q(N206)
         );
  DFQRM1SA add_regs_reg_8__8_ ( .D(intadd_7_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[72]) );
  DFQRM1SA add_regs_reg_8__7_ ( .D(N80), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[71]) );
  DFQRM1SA add_regs_reg_8__6_ ( .D(N79), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[70]) );
  DFQRM1SA add_regs_reg_8__5_ ( .D(N78), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[69]) );
  DFQRM1SA add_regs_reg_8__3_ ( .D(N76), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[67]) );
  DFQRM1SA add_regs_reg_8__2_ ( .D(N75), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[66]) );
  DFQRM1SA add_regs_reg_8__1_ ( .D(N74), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[65]) );
  DFQRM1SA add_regs_reg_8__0_ ( .D(N73), .CK(CLK_Filter), .RB(rst_n), .Q(N189)
         );
  DFQRM1SA add_regs_reg_7__8_ ( .D(intadd_8_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[64]) );
  DFQRM1SA add_regs_reg_7__7_ ( .D(N71), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[63]) );
  DFQRM1SA add_regs_reg_7__6_ ( .D(N70), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[62]) );
  DFQRM1SA add_regs_reg_7__5_ ( .D(N69), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[61]) );
  DFQRM1SA add_regs_reg_7__4_ ( .D(N68), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[60]) );
  DFQRM1SA add_regs_reg_7__3_ ( .D(N67), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[59]) );
  DFQRM1SA add_regs_reg_7__2_ ( .D(N66), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[58]) );
  DFQRM1SA add_regs_reg_7__1_ ( .D(N65), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[57]) );
  DFQRM1SA add_regs_reg_7__0_ ( .D(N64), .CK(CLK_Filter), .RB(rst_n), .Q(N173)
         );
  DFQRM1SA add_regs_reg_6__8_ ( .D(intadd_9_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[56]) );
  DFQRM1SA add_regs_reg_6__6_ ( .D(N61), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[54]) );
  DFQRM1SA add_regs_reg_6__5_ ( .D(N60), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[53]) );
  DFQRM1SA add_regs_reg_6__4_ ( .D(N59), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[52]) );
  DFQRM1SA add_regs_reg_6__3_ ( .D(N58), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[51]) );
  DFQRM1SA add_regs_reg_6__2_ ( .D(N57), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[50]) );
  DFQRM1SA add_regs_reg_6__1_ ( .D(N56), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[49]) );
  DFQRM1SA add_regs_reg_6__0_ ( .D(N55), .CK(CLK_Filter), .RB(rst_n), .Q(N158)
         );
  DFQRM1SA add_regs_reg_5__8_ ( .D(intadd_10_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[48]) );
  DFQRM1SA add_regs_reg_5__7_ ( .D(N53), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[47]) );
  DFQRM1SA add_regs_reg_5__6_ ( .D(N52), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[46]) );
  DFQRM1SA add_regs_reg_5__5_ ( .D(N51), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[45]) );
  DFQRM1SA add_regs_reg_5__4_ ( .D(N50), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[44]) );
  DFQRM1SA add_regs_reg_5__3_ ( .D(N49), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[43]) );
  DFQRM1SA add_regs_reg_5__2_ ( .D(N48), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[42]) );
  DFQRM1SA add_regs_reg_5__0_ ( .D(N46), .CK(CLK_Filter), .RB(rst_n), .Q(N144)
         );
  DFQRM1SA add_regs_reg_4__8_ ( .D(intadd_11_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[40]) );
  DFQRM1SA add_regs_reg_4__7_ ( .D(N44), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[39]) );
  DFQRM1SA add_regs_reg_4__6_ ( .D(N43), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[38]) );
  DFQRM1SA add_regs_reg_4__5_ ( .D(N42), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[37]) );
  DFQRM1SA add_regs_reg_4__4_ ( .D(N41), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[36]) );
  DFQRM1SA add_regs_reg_4__3_ ( .D(N40), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[35]) );
  DFQRM1SA add_regs_reg_4__2_ ( .D(N39), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[34]) );
  DFQRM1SA add_regs_reg_4__1_ ( .D(N38), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[33]) );
  DFQRM1SA add_regs_reg_4__0_ ( .D(N37), .CK(CLK_Filter), .RB(rst_n), .Q(N127)
         );
  DFQRM1SA add_regs_reg_3__8_ ( .D(intadd_12_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[32]) );
  DFQRM1SA add_regs_reg_3__7_ ( .D(N35), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[31]) );
  DFQRM1SA add_regs_reg_3__6_ ( .D(N34), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[30]) );
  DFQRM1SA add_regs_reg_3__5_ ( .D(N33), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[29]) );
  DFQRM1SA add_regs_reg_3__3_ ( .D(N31), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[27]) );
  DFQRM1SA add_regs_reg_3__2_ ( .D(N30), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[26]) );
  DFQRM1SA add_regs_reg_3__1_ ( .D(N29), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[25]) );
  DFQRM1SA add_regs_reg_3__0_ ( .D(N28), .CK(CLK_Filter), .RB(rst_n), .Q(N115)
         );
  DFQRM1SA add_regs_reg_2__8_ ( .D(intadd_13_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[24]) );
  DFQRM1SA add_regs_reg_2__7_ ( .D(N26), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[23]) );
  DFQRM1SA add_regs_reg_2__6_ ( .D(N25), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[22]) );
  DFQRM1SA add_regs_reg_2__5_ ( .D(N24), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[21]) );
  DFQRM1SA add_regs_reg_2__4_ ( .D(N23), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[20]) );
  DFQRM1SA add_regs_reg_2__2_ ( .D(N21), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[18]) );
  DFQRM1SA add_regs_reg_2__1_ ( .D(N20), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[17]) );
  DFQRM1SA add_regs_reg_2__0_ ( .D(N19), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[16]) );
  DFQRM1SA add_regs_reg_1__8_ ( .D(intadd_14_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[15]) );
  DFQRM1SA add_regs_reg_1__7_ ( .D(N17), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[14]) );
  DFQRM1SA add_regs_reg_1__6_ ( .D(N16), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[13]) );
  DFQRM1SA add_regs_reg_1__5_ ( .D(N15), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[12]) );
  DFQRM1SA add_regs_reg_1__4_ ( .D(N14), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[11]) );
  DFQRM1SA add_regs_reg_1__3_ ( .D(N13), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[10]) );
  DFQRM1SA add_regs_reg_1__2_ ( .D(N12), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[9]) );
  DFQRM1SA add_regs_reg_1__0_ ( .D(N10), .CK(CLK_Filter), .RB(rst_n), .Q(N101)
         );
  DFQRM1SA add_regs_reg_0__8_ ( .D(intadd_15_n1), .CK(CLK_Filter), .RB(rst_n), 
        .Q(add_regs[8]) );
  DFQRM1SA add_regs_reg_0__7_ ( .D(N8), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[7]) );
  DFQRM1SA add_regs_reg_0__6_ ( .D(N7), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[6]) );
  DFQRM1SA add_regs_reg_0__5_ ( .D(N6), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[5]) );
  DFQRM1SA add_regs_reg_0__4_ ( .D(N5), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[4]) );
  DFQRM1SA add_regs_reg_0__3_ ( .D(N4), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[3]) );
  DFQRM1SA add_regs_reg_0__2_ ( .D(N3), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[2]) );
  DFQRM1SA add_regs_reg_0__1_ ( .D(N2), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[1]) );
  DFQRM1SA add_regs_reg_0__0_ ( .D(N1), .CK(CLK_Filter), .RB(rst_n), .Q(
        add_regs[0]) );
  ADFM1SA intadd_0_U2 ( .A(intadd_0_A_17_), .B(intadd_26_n1), .CI(intadd_0_n2), 
        .CO(intadd_0_n1), .S(N415) );
  ADFM1SA intadd_0_U3 ( .A(intadd_0_A_16_), .B(intadd_27_n1), .CI(intadd_0_n3), 
        .CO(intadd_0_n2), .S(N414) );
  ADFM1SA intadd_0_U4 ( .A(intadd_0_A_15_), .B(intadd_17_n1), .CI(intadd_0_n4), 
        .CO(intadd_0_n3), .S(N413) );
  ADFM1SA intadd_0_U5 ( .A(intadd_0_A_14_), .B(intadd_18_n1), .CI(intadd_0_n5), 
        .CO(intadd_0_n4), .S(N412) );
  ADFM1SA intadd_0_U6 ( .A(intadd_0_A_13_), .B(intadd_19_n1), .CI(intadd_0_n6), 
        .CO(intadd_0_n5), .S(N411) );
  ADFM1SA intadd_0_U7 ( .A(intadd_0_A_12_), .B(intadd_20_n1), .CI(intadd_0_n7), 
        .CO(intadd_0_n6), .S(N410) );
  ADFM1SA intadd_0_U8 ( .A(intadd_0_A_11_), .B(intadd_21_n1), .CI(intadd_0_n8), 
        .CO(intadd_0_n7), .S(N409) );
  ADFM1SA intadd_0_U9 ( .A(intadd_0_A_10_), .B(intadd_22_n1), .CI(intadd_0_n9), 
        .CO(intadd_0_n8), .S(N408) );
  ADFM1SA intadd_0_U10 ( .A(intadd_0_A_9_), .B(intadd_23_n1), .CI(intadd_0_n10), .CO(intadd_0_n9), .S(N407) );
  ADFM1SA intadd_0_U11 ( .A(intadd_0_A_8_), .B(intadd_24_n1), .CI(intadd_0_n11), .CO(intadd_0_n10), .S(N406) );
  ADFM1SA intadd_0_U12 ( .A(intadd_0_A_7_), .B(intadd_28_n1), .CI(intadd_0_n12), .CO(intadd_0_n11), .S(N405) );
  ADFM1SA intadd_0_U13 ( .A(intadd_0_A_6_), .B(intadd_29_n1), .CI(intadd_0_n13), .CO(intadd_0_n12), .S(N404) );
  ADFM1SA intadd_0_U14 ( .A(intadd_0_A_5_), .B(intadd_0_B_5_), .CI(
        intadd_0_n14), .CO(intadd_0_n13), .S(N403) );
  ADFM1SA intadd_0_U16 ( .A(intadd_0_A_3_), .B(intadd_0_B_3_), .CI(
        intadd_0_n16), .CO(intadd_0_n15), .S(N401) );
  ADFM1SA intadd_0_U17 ( .A(intadd_0_A_2_), .B(intadd_0_B_2_), .CI(
        intadd_0_n17), .CO(intadd_0_n16), .S(N400) );
  ADFM1SA intadd_0_U18 ( .A(intadd_0_A_1_), .B(intadd_0_B_1_), .CI(
        intadd_0_n18), .CO(intadd_0_n17), .S(N399) );
  ADFM1SA intadd_0_U19 ( .A(order[101]), .B(order[42]), .CI(order[85]), .CO(
        intadd_0_n18), .S(N398) );
  ADFM1SA intadd_4_U2 ( .A(intadd_4_A_6_), .B(intadd_4_B_6_), .CI(intadd_4_n2), 
        .CO(intadd_4_n1), .S(N185) );
  ADFM1SA intadd_4_U3 ( .A(intadd_4_A_5_), .B(intadd_4_B_5_), .CI(intadd_4_n3), 
        .CO(intadd_4_n2), .S(N184) );
  ADFM1SA intadd_4_U4 ( .A(intadd_4_A_4_), .B(intadd_4_B_4_), .CI(intadd_4_n4), 
        .CO(intadd_4_n3), .S(N183) );
  ADFM1SA intadd_4_U5 ( .A(intadd_4_A_3_), .B(intadd_4_B_3_), .CI(intadd_4_n5), 
        .CO(intadd_4_n4), .S(N182) );
  ADFM1SA intadd_4_U6 ( .A(intadd_4_A_2_), .B(intadd_4_B_2_), .CI(intadd_4_n6), 
        .CO(intadd_4_n5), .S(N181) );
  ADFM1SA intadd_4_U7 ( .A(intadd_4_A_1_), .B(intadd_4_B_1_), .CI(intadd_4_n7), 
        .CO(intadd_4_n6), .S(N180) );
  ADFM1SA intadd_31_U2 ( .A(intadd_31_A_3_), .B(intadd_31_B_3_), .CI(
        intadd_31_n2), .CO(intadd_31_n1), .S(N168) );
  ADFM1SA intadd_31_U3 ( .A(intadd_31_A_2_), .B(intadd_31_B_2_), .CI(
        intadd_31_n3), .CO(intadd_31_n2), .S(N167) );
  ADFM1SA intadd_31_U4 ( .A(intadd_31_A_1_), .B(intadd_31_B_1_), .CI(
        intadd_31_n4), .CO(intadd_31_n3), .S(N166) );
  ADFM1SA intadd_1_U2 ( .A(add_regs[39]), .B(intadd_1_B_9_), .CI(intadd_1_n2), 
        .CO(intadd_1_n1), .S(N139) );
  ADFM1SA intadd_1_U3 ( .A(intadd_1_A_8_), .B(intadd_1_B_8_), .CI(intadd_1_n3), 
        .CO(intadd_1_n2), .S(N138) );
  ADFM1SA intadd_1_U4 ( .A(intadd_1_A_7_), .B(intadd_1_B_7_), .CI(intadd_1_n4), 
        .CO(intadd_1_n3), .S(N137) );
  ADFM1SA intadd_1_U5 ( .A(intadd_1_A_6_), .B(intadd_1_B_6_), .CI(intadd_1_n5), 
        .CO(intadd_1_n4), .S(N136) );
  ADFM1SA intadd_1_U6 ( .A(intadd_1_A_5_), .B(intadd_1_B_5_), .CI(intadd_1_n6), 
        .CO(intadd_1_n5), .S(N135) );
  ADFM1SA intadd_1_U7 ( .A(intadd_1_A_4_), .B(intadd_1_B_4_), .CI(intadd_1_n7), 
        .CO(intadd_1_n6), .S(N134) );
  ADFM1SA intadd_1_U8 ( .A(intadd_1_A_3_), .B(intadd_1_B_3_), .CI(intadd_1_n8), 
        .CO(intadd_1_n7), .S(N133) );
  ADFM1SA intadd_1_U9 ( .A(intadd_1_A_2_), .B(intadd_1_B_2_), .CI(intadd_1_n9), 
        .CO(intadd_1_n8), .S(N132) );
  ADFM1SA intadd_1_U11 ( .A(N127), .B(intadd_1_B_0_), .CI(intadd_1_CI), .CO(
        intadd_1_n10), .S(N130) );
  ADFM1SA intadd_16_U2 ( .A(add_regs[13]), .B(add_regs[15]), .CI(intadd_16_n2), 
        .CO(intadd_16_n1), .S(N109) );
  ADFM1SA intadd_16_U3 ( .A(add_regs[12]), .B(add_regs[14]), .CI(intadd_16_n3), 
        .CO(intadd_16_n2), .S(N108) );
  ADFM1SA intadd_16_U4 ( .A(add_regs[11]), .B(add_regs[13]), .CI(intadd_16_n4), 
        .CO(intadd_16_n3), .S(N107) );
  ADFM1SA intadd_16_U5 ( .A(add_regs[10]), .B(add_regs[12]), .CI(intadd_16_n5), 
        .CO(intadd_16_n4), .S(N106) );
  ADFM1SA intadd_16_U6 ( .A(add_regs[9]), .B(add_regs[11]), .CI(intadd_16_n6), 
        .CO(intadd_16_n5), .S(N105) );
  ADFM1SA intadd_16_U7 ( .A(N102), .B(add_regs[10]), .CI(intadd_16_CI), .CO(
        intadd_16_n6), .S(N104) );
  ADFM1SA intadd_5_U2 ( .A(shift_regs[95]), .B(shift_regs[87]), .CI(
        intadd_5_n2), .CO(intadd_5_n1), .S(N98) );
  ADFM1SA intadd_5_U3 ( .A(shift_regs[94]), .B(shift_regs[86]), .CI(
        intadd_5_n3), .CO(intadd_5_n2), .S(N97) );
  ADFM1SA intadd_5_U4 ( .A(shift_regs[93]), .B(shift_regs[85]), .CI(
        intadd_5_n4), .CO(intadd_5_n3), .S(N96) );
  ADFM1SA intadd_5_U5 ( .A(shift_regs[92]), .B(shift_regs[84]), .CI(
        intadd_5_n5), .CO(intadd_5_n4), .S(N95) );
  ADFM1SA intadd_5_U6 ( .A(shift_regs[91]), .B(shift_regs[83]), .CI(
        intadd_5_n6), .CO(intadd_5_n5), .S(N94) );
  ADFM1SA intadd_5_U7 ( .A(shift_regs[90]), .B(shift_regs[82]), .CI(
        intadd_5_n7), .CO(intadd_5_n6), .S(N93) );
  ADFM1SA intadd_5_U8 ( .A(shift_regs[89]), .B(shift_regs[81]), .CI(
        intadd_5_CI), .CO(intadd_5_n7), .S(N92) );
  ADFM1SA intadd_6_U2 ( .A(shift_regs[103]), .B(shift_regs[79]), .CI(
        intadd_6_n2), .CO(intadd_6_n1), .S(N89) );
  ADFM1SA intadd_6_U3 ( .A(shift_regs[102]), .B(shift_regs[78]), .CI(
        intadd_6_n3), .CO(intadd_6_n2), .S(N88) );
  ADFM1SA intadd_6_U4 ( .A(shift_regs[101]), .B(shift_regs[77]), .CI(
        intadd_6_n4), .CO(intadd_6_n3), .S(N87) );
  ADFM1SA intadd_6_U5 ( .A(shift_regs[100]), .B(shift_regs[76]), .CI(
        intadd_6_n5), .CO(intadd_6_n4), .S(N86) );
  ADFM1SA intadd_6_U6 ( .A(shift_regs[99]), .B(shift_regs[75]), .CI(
        intadd_6_n6), .CO(intadd_6_n5), .S(N85) );
  ADFM1SA intadd_6_U7 ( .A(shift_regs[98]), .B(shift_regs[74]), .CI(
        intadd_6_n7), .CO(intadd_6_n6), .S(N84) );
  ADFM1SA intadd_6_U8 ( .A(shift_regs[97]), .B(shift_regs[73]), .CI(
        intadd_6_CI), .CO(intadd_6_n7), .S(N83) );
  ADFM1SA intadd_7_U2 ( .A(shift_regs[111]), .B(shift_regs[71]), .CI(
        intadd_7_n2), .CO(intadd_7_n1), .S(N80) );
  ADFM1SA intadd_7_U3 ( .A(shift_regs[110]), .B(shift_regs[70]), .CI(
        intadd_7_n3), .CO(intadd_7_n2), .S(N79) );
  ADFM1SA intadd_7_U4 ( .A(shift_regs[109]), .B(shift_regs[69]), .CI(
        intadd_7_n4), .CO(intadd_7_n3), .S(N78) );
  ADFM1SA intadd_7_U6 ( .A(shift_regs[107]), .B(shift_regs[67]), .CI(
        intadd_7_n6), .CO(intadd_7_n5), .S(N76) );
  ADFM1SA intadd_7_U7 ( .A(shift_regs[106]), .B(shift_regs[66]), .CI(
        intadd_7_n7), .CO(intadd_7_n6), .S(N75) );
  ADFM1SA intadd_7_U8 ( .A(shift_regs[105]), .B(shift_regs[65]), .CI(
        intadd_7_CI), .CO(intadd_7_n7), .S(N74) );
  ADFM1SA intadd_8_U2 ( .A(shift_regs[119]), .B(shift_regs[63]), .CI(
        intadd_8_n2), .CO(intadd_8_n1), .S(N71) );
  ADFM1SA intadd_8_U3 ( .A(shift_regs[118]), .B(shift_regs[62]), .CI(
        intadd_8_n3), .CO(intadd_8_n2), .S(N70) );
  ADFM1SA intadd_8_U4 ( .A(shift_regs[117]), .B(shift_regs[61]), .CI(
        intadd_8_n4), .CO(intadd_8_n3), .S(N69) );
  ADFM1SA intadd_8_U5 ( .A(shift_regs[116]), .B(shift_regs[60]), .CI(
        intadd_8_n5), .CO(intadd_8_n4), .S(N68) );
  ADFM1SA intadd_8_U6 ( .A(shift_regs[115]), .B(shift_regs[59]), .CI(
        intadd_8_n6), .CO(intadd_8_n5), .S(N67) );
  ADFM1SA intadd_8_U7 ( .A(shift_regs[114]), .B(shift_regs[58]), .CI(
        intadd_8_n7), .CO(intadd_8_n6), .S(N66) );
  ADFM1SA intadd_8_U8 ( .A(shift_regs[113]), .B(shift_regs[57]), .CI(
        intadd_8_CI), .CO(intadd_8_n7), .S(N65) );
  ADFM1SA intadd_9_U2 ( .A(shift_regs[127]), .B(shift_regs[55]), .CI(
        intadd_9_n2), .CO(intadd_9_n1), .S(N62) );
  ADFM1SA intadd_9_U3 ( .A(shift_regs[126]), .B(shift_regs[54]), .CI(
        intadd_9_n3), .CO(intadd_9_n2), .S(N61) );
  ADFM1SA intadd_9_U4 ( .A(shift_regs[125]), .B(shift_regs[53]), .CI(
        intadd_9_n4), .CO(intadd_9_n3), .S(N60) );
  ADFM1SA intadd_9_U5 ( .A(shift_regs[124]), .B(shift_regs[52]), .CI(
        intadd_9_n5), .CO(intadd_9_n4), .S(N59) );
  ADFM1SA intadd_9_U6 ( .A(shift_regs[123]), .B(shift_regs[51]), .CI(
        intadd_9_n6), .CO(intadd_9_n5), .S(N58) );
  ADFM1SA intadd_9_U7 ( .A(shift_regs[122]), .B(shift_regs[50]), .CI(
        intadd_9_n7), .CO(intadd_9_n6), .S(N57) );
  ADFM1SA intadd_9_U8 ( .A(shift_regs[121]), .B(shift_regs[49]), .CI(
        intadd_9_CI), .CO(intadd_9_n7), .S(N56) );
  ADFM1SA intadd_10_U2 ( .A(shift_regs[135]), .B(shift_regs[47]), .CI(
        intadd_10_n2), .CO(intadd_10_n1), .S(N53) );
  ADFM1SA intadd_10_U3 ( .A(shift_regs[134]), .B(shift_regs[46]), .CI(
        intadd_10_n3), .CO(intadd_10_n2), .S(N52) );
  ADFM1SA intadd_10_U4 ( .A(shift_regs[133]), .B(shift_regs[45]), .CI(
        intadd_10_n4), .CO(intadd_10_n3), .S(N51) );
  ADFM1SA intadd_10_U5 ( .A(shift_regs[132]), .B(shift_regs[44]), .CI(
        intadd_10_n5), .CO(intadd_10_n4), .S(N50) );
  ADFM1SA intadd_10_U6 ( .A(shift_regs[131]), .B(shift_regs[43]), .CI(
        intadd_10_n6), .CO(intadd_10_n5), .S(N49) );
  ADFM1SA intadd_10_U7 ( .A(shift_regs[130]), .B(shift_regs[42]), .CI(
        intadd_10_n7), .CO(intadd_10_n6), .S(N48) );
  ADFM1SA intadd_11_U2 ( .A(shift_regs[143]), .B(shift_regs[39]), .CI(
        intadd_11_n2), .CO(intadd_11_n1), .S(N44) );
  ADFM1SA intadd_11_U3 ( .A(shift_regs[142]), .B(shift_regs[38]), .CI(
        intadd_11_n3), .CO(intadd_11_n2), .S(N43) );
  ADFM1SA intadd_11_U4 ( .A(shift_regs[141]), .B(shift_regs[37]), .CI(
        intadd_11_n4), .CO(intadd_11_n3), .S(N42) );
  ADFM1SA intadd_11_U5 ( .A(shift_regs[140]), .B(shift_regs[36]), .CI(
        intadd_11_n5), .CO(intadd_11_n4), .S(N41) );
  ADFM1SA intadd_11_U6 ( .A(shift_regs[139]), .B(shift_regs[35]), .CI(
        intadd_11_n6), .CO(intadd_11_n5), .S(N40) );
  ADFM1SA intadd_11_U7 ( .A(shift_regs[138]), .B(shift_regs[34]), .CI(
        intadd_11_n7), .CO(intadd_11_n6), .S(N39) );
  ADFM1SA intadd_11_U8 ( .A(shift_regs[137]), .B(shift_regs[33]), .CI(
        intadd_11_CI), .CO(intadd_11_n7), .S(N38) );
  ADFM1SA intadd_12_U2 ( .A(shift_regs[151]), .B(shift_regs[31]), .CI(
        intadd_12_n2), .CO(intadd_12_n1), .S(N35) );
  ADFM1SA intadd_12_U3 ( .A(shift_regs[150]), .B(shift_regs[30]), .CI(
        intadd_12_n3), .CO(intadd_12_n2), .S(N34) );
  ADFM1SA intadd_12_U4 ( .A(shift_regs[149]), .B(shift_regs[29]), .CI(
        intadd_12_n4), .CO(intadd_12_n3), .S(N33) );
  ADFM1SA intadd_12_U6 ( .A(shift_regs[147]), .B(shift_regs[27]), .CI(
        intadd_12_n6), .CO(intadd_12_n5), .S(N31) );
  ADFM1SA intadd_12_U7 ( .A(shift_regs[146]), .B(shift_regs[26]), .CI(
        intadd_12_n7), .CO(intadd_12_n6), .S(N30) );
  ADFM1SA intadd_12_U8 ( .A(shift_regs[145]), .B(shift_regs[25]), .CI(
        intadd_12_CI), .CO(intadd_12_n7), .S(N29) );
  ADFM1SA intadd_13_U2 ( .A(shift_regs[159]), .B(shift_regs[23]), .CI(
        intadd_13_n2), .CO(intadd_13_n1), .S(N26) );
  ADFM1SA intadd_13_U3 ( .A(shift_regs[158]), .B(shift_regs[22]), .CI(
        intadd_13_n3), .CO(intadd_13_n2), .S(N25) );
  ADFM1SA intadd_13_U4 ( .A(shift_regs[157]), .B(shift_regs[21]), .CI(
        intadd_13_n4), .CO(intadd_13_n3), .S(N24) );
  ADFM1SA intadd_13_U5 ( .A(shift_regs[156]), .B(shift_regs[20]), .CI(
        intadd_13_n5), .CO(intadd_13_n4), .S(N23) );
  ADFM1SA intadd_13_U7 ( .A(shift_regs[154]), .B(shift_regs[18]), .CI(
        intadd_13_n7), .CO(intadd_13_n6), .S(N21) );
  ADFM1SA intadd_13_U8 ( .A(shift_regs[153]), .B(shift_regs[17]), .CI(
        intadd_13_CI), .CO(intadd_13_n7), .S(N20) );
  ADFM1SA intadd_14_U2 ( .A(shift_regs[167]), .B(shift_regs[15]), .CI(
        intadd_14_n2), .CO(intadd_14_n1), .S(N17) );
  ADFM1SA intadd_14_U3 ( .A(shift_regs[166]), .B(shift_regs[14]), .CI(
        intadd_14_n3), .CO(intadd_14_n2), .S(N16) );
  ADFM1SA intadd_14_U4 ( .A(shift_regs[165]), .B(shift_regs[13]), .CI(
        intadd_14_n4), .CO(intadd_14_n3), .S(N15) );
  ADFM1SA intadd_14_U5 ( .A(shift_regs[164]), .B(shift_regs[12]), .CI(
        intadd_14_n5), .CO(intadd_14_n4), .S(N14) );
  ADFM1SA intadd_14_U6 ( .A(shift_regs[163]), .B(shift_regs[11]), .CI(
        intadd_14_n6), .CO(intadd_14_n5), .S(N13) );
  ADFM1SA intadd_14_U7 ( .A(shift_regs[162]), .B(shift_regs[10]), .CI(
        intadd_14_n7), .CO(intadd_14_n6), .S(N12) );
  ADFM1SA intadd_15_U2 ( .A(shift_regs[175]), .B(shift_regs[7]), .CI(
        intadd_15_n2), .CO(intadd_15_n1), .S(N8) );
  ADFM1SA intadd_15_U3 ( .A(shift_regs[174]), .B(shift_regs[6]), .CI(
        intadd_15_n3), .CO(intadd_15_n2), .S(N7) );
  ADFM1SA intadd_15_U4 ( .A(shift_regs[173]), .B(shift_regs[5]), .CI(
        intadd_15_n4), .CO(intadd_15_n3), .S(N6) );
  ADFM1SA intadd_15_U5 ( .A(shift_regs[172]), .B(shift_regs[4]), .CI(
        intadd_15_n5), .CO(intadd_15_n4), .S(N5) );
  ADFM1SA intadd_15_U6 ( .A(shift_regs[171]), .B(shift_regs[3]), .CI(
        intadd_15_n6), .CO(intadd_15_n5), .S(N4) );
  ADFM1SA intadd_15_U7 ( .A(shift_regs[170]), .B(shift_regs[2]), .CI(
        intadd_15_n7), .CO(intadd_15_n6), .S(N3) );
  ADFM1SA intadd_15_U8 ( .A(shift_regs[169]), .B(shift_regs[1]), .CI(
        intadd_15_CI), .CO(intadd_15_n7), .S(N2) );
  ADFM1SA intadd_0_U15 ( .A(intadd_0_A_4_), .B(intadd_35_n1), .CI(intadd_0_n15), .CO(intadd_0_n14), .S(N402) );
  ADFM1SA intadd_4_U8 ( .A(N173), .B(intadd_4_B_0_), .CI(intadd_4_CI), .CO(
        intadd_4_n7), .S(N179) );
  ADFM1SA intadd_1_U10 ( .A(intadd_1_A_1_), .B(intadd_1_B_1_), .CI(
        intadd_1_n10), .CO(intadd_1_n9), .S(N131) );
  ADFM1SA intadd_7_U5 ( .A(shift_regs[108]), .B(shift_regs[68]), .CI(
        intadd_7_n5), .CO(intadd_7_n4), .S(N77) );
  ADFM1SA intadd_10_U8 ( .A(shift_regs[129]), .B(shift_regs[41]), .CI(
        intadd_10_CI), .CO(intadd_10_n7), .S(N47) );
  ADFM1SA intadd_12_U5 ( .A(shift_regs[148]), .B(shift_regs[28]), .CI(
        intadd_12_n5), .CO(intadd_12_n4), .S(N32) );
  ADFM1SA intadd_13_U6 ( .A(shift_regs[155]), .B(shift_regs[19]), .CI(
        intadd_13_n6), .CO(intadd_13_n5), .S(N22) );
  ADFM1SA intadd_14_U8 ( .A(shift_regs[161]), .B(shift_regs[9]), .CI(
        intadd_14_CI), .CO(intadd_14_n7), .S(N11) );
  ADFM1SA intadd_26_U2 ( .A(intadd_26_A_3_), .B(intadd_26_B_3_), .CI(
        intadd_26_n2), .CO(intadd_26_n1), .S(intadd_0_A_16_) );
  ADFM1SA intadd_27_U2 ( .A(intadd_26_SUM_2_), .B(intadd_27_B_3_), .CI(
        intadd_27_n2), .CO(intadd_27_n1), .S(intadd_0_A_15_) );
  ADFM1SA intadd_17_U2 ( .A(intadd_17_A_4_), .B(intadd_34_n1), .CI(
        intadd_17_n2), .CO(intadd_17_n1), .S(intadd_0_A_14_) );
  ADFM1SA intadd_18_U2 ( .A(intadd_18_A_4_), .B(intadd_17_SUM_3_), .CI(
        intadd_18_n2), .CO(intadd_18_n1), .S(intadd_0_A_13_) );
  ADFM1SA intadd_19_U2 ( .A(intadd_18_SUM_3_), .B(intadd_17_SUM_2_), .CI(
        intadd_19_n2), .CO(intadd_19_n1), .S(intadd_0_A_12_) );
  ADFM1SA intadd_20_U2 ( .A(intadd_19_SUM_3_), .B(intadd_18_SUM_2_), .CI(
        intadd_20_n2), .CO(intadd_20_n1), .S(intadd_0_A_11_) );
  ADFM1SA intadd_21_U2 ( .A(intadd_20_SUM_3_), .B(intadd_19_SUM_2_), .CI(
        intadd_21_n2), .CO(intadd_21_n1), .S(intadd_0_A_10_) );
  ADFM1SA intadd_22_U2 ( .A(intadd_21_SUM_3_), .B(intadd_20_SUM_2_), .CI(
        intadd_22_n2), .CO(intadd_22_n1), .S(intadd_0_A_9_) );
  ADFM1SA intadd_23_U2 ( .A(intadd_22_SUM_3_), .B(intadd_21_SUM_2_), .CI(
        intadd_23_n2), .CO(intadd_23_n1), .S(intadd_0_A_8_) );
  ADFM1SA intadd_24_U2 ( .A(intadd_23_SUM_3_), .B(intadd_22_SUM_2_), .CI(
        intadd_24_n2), .CO(intadd_24_n1), .S(intadd_0_A_7_) );
  ADFM1SA intadd_28_U2 ( .A(intadd_24_SUM_3_), .B(intadd_23_SUM_2_), .CI(
        intadd_28_n2), .CO(intadd_28_n1), .S(intadd_0_A_6_) );
  ADFM1SA intadd_29_U2 ( .A(intadd_28_SUM_2_), .B(intadd_24_SUM_2_), .CI(
        intadd_29_n2), .CO(intadd_29_n1), .S(intadd_0_A_5_) );
  ADFM1SA intadd_35_U2 ( .A(intadd_29_SUM_1_), .B(intadd_35_B_2_), .CI(
        intadd_35_n2), .CO(intadd_35_n1), .S(intadd_0_A_3_) );
  ADFM1SA intadd_35_U3 ( .A(intadd_35_A_1_), .B(intadd_35_B_1_), .CI(
        intadd_35_n3), .CO(intadd_35_n2), .S(intadd_0_B_2_) );
  ADFM1SA intadd_35_U4 ( .A(order[9]), .B(order[0]), .CI(order[102]), .CO(
        intadd_35_n3), .S(intadd_0_B_1_) );
  DFQRM1SA order_reg_8__0_ ( .D(N189), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[101]) );
  DFQRM1SA order_reg_4__0_ ( .D(N127), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[42]) );
  DFQRM1SA order_reg_7__0_ ( .D(N173), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[85]) );
  ADFM1SA intadd_2_U2 ( .A(intadd_2_A_7_), .B(intadd_2_B_7_), .CI(intadd_2_n2), 
        .CO(intadd_2_n1), .S(intadd_2_SUM_7_) );
  ADFM1SA intadd_2_U3 ( .A(intadd_2_A_6_), .B(intadd_2_B_6_), .CI(intadd_2_n3), 
        .CO(intadd_2_n2), .S(intadd_2_SUM_6_) );
  ADFM1SA intadd_2_U4 ( .A(intadd_2_A_5_), .B(intadd_2_B_5_), .CI(intadd_2_n4), 
        .CO(intadd_2_n3), .S(intadd_2_SUM_5_) );
  ADFM1SA intadd_2_U5 ( .A(intadd_2_A_4_), .B(intadd_2_B_4_), .CI(intadd_2_n5), 
        .CO(intadd_2_n4), .S(intadd_2_SUM_4_) );
  ADFM1SA intadd_2_U6 ( .A(intadd_2_A_3_), .B(intadd_2_B_3_), .CI(intadd_2_n6), 
        .CO(intadd_2_n5), .S(intadd_2_SUM_3_) );
  ADFM1SA intadd_2_U7 ( .A(add_regs[74]), .B(intadd_2_B_2_), .CI(intadd_2_n7), 
        .CO(intadd_2_n6), .S(intadd_2_SUM_2_) );
  ADFM1SA intadd_2_U9 ( .A(N207), .B(intadd_2_B_0_), .CI(intadd_2_CI), .CO(
        intadd_2_n8), .S(intadd_2_SUM_0_) );
  ADFM1SA intadd_3_U2 ( .A(intadd_3_A_6_), .B(intadd_3_B_6_), .CI(intadd_3_n2), 
        .CO(intadd_3_n1), .S(intadd_3_SUM_6_) );
  ADFM1SA intadd_3_U3 ( .A(intadd_3_A_5_), .B(intadd_3_B_5_), .CI(intadd_3_n3), 
        .CO(intadd_3_n2), .S(intadd_3_SUM_5_) );
  ADFM1SA intadd_3_U4 ( .A(intadd_3_A_4_), .B(intadd_3_B_4_), .CI(intadd_3_n4), 
        .CO(intadd_3_n3), .S(intadd_3_SUM_4_) );
  ADFM1SA intadd_3_U5 ( .A(intadd_3_A_3_), .B(intadd_3_B_3_), .CI(intadd_3_n5), 
        .CO(intadd_3_n4), .S(intadd_3_SUM_3_) );
  ADFM1SA intadd_3_U6 ( .A(intadd_3_A_2_), .B(intadd_3_B_2_), .CI(intadd_3_n6), 
        .CO(intadd_3_n5), .S(intadd_3_SUM_2_) );
  ADFM1SA intadd_3_U7 ( .A(intadd_3_A_1_), .B(intadd_3_B_1_), .CI(intadd_3_n7), 
        .CO(intadd_3_n6), .S(intadd_3_SUM_1_) );
  ADFM1SA intadd_32_U2 ( .A(intadd_32_A_3_), .B(intadd_32_B_3_), .CI(
        intadd_32_n2), .CO(intadd_32_n1), .S(intadd_32_SUM_3_) );
  ADFM1SA intadd_31_U5 ( .A(add_regs[50]), .B(add_regs[52]), .CI(intadd_31_CI), 
        .CO(intadd_31_n4), .S(intadd_31_SUM_0_) );
  ADFM1SA intadd_32_U4 ( .A(intadd_32_A_1_), .B(intadd_32_B_1_), .CI(
        intadd_32_n4), .CO(intadd_32_n3), .S(intadd_32_SUM_1_) );
  ADFM1SA intadd_32_U5 ( .A(add_regs[52]), .B(intadd_32_B_0_), .CI(
        intadd_32_CI), .CO(intadd_32_n4), .S(intadd_32_SUM_0_) );
  ADFM1SA intadd_30_U2 ( .A(add_regs[48]), .B(intadd_30_B_3_), .CI(
        intadd_30_n2), .CO(intadd_30_n1), .S(intadd_30_SUM_3_) );
  ADFM1SA intadd_30_U3 ( .A(add_regs[47]), .B(intadd_30_B_2_), .CI(
        intadd_30_n3), .CO(intadd_30_n2), .S(intadd_30_SUM_2_) );
  ADFM1SA intadd_30_U4 ( .A(add_regs[46]), .B(intadd_30_B_1_), .CI(
        intadd_30_n4), .CO(intadd_30_n3), .S(intadd_30_SUM_1_) );
  ADFM1SA intadd_30_U5 ( .A(add_regs[45]), .B(intadd_30_B_0_), .CI(
        intadd_30_CI), .CO(intadd_30_n4), .S(intadd_30_SUM_0_) );
  ADFM1SA intadd_25_U2 ( .A(add_regs[32]), .B(intadd_25_B_4_), .CI(
        intadd_25_n2), .CO(intadd_25_n1), .S(intadd_25_SUM_4_) );
  ADFM1SA intadd_25_U3 ( .A(add_regs[31]), .B(intadd_25_B_3_), .CI(
        intadd_25_n3), .CO(intadd_25_n2), .S(intadd_25_SUM_3_) );
  ADFM1SA intadd_25_U4 ( .A(add_regs[30]), .B(intadd_25_B_2_), .CI(
        intadd_25_n4), .CO(intadd_25_n3), .S(intadd_25_SUM_2_) );
  ADFM1SA intadd_25_U5 ( .A(intadd_25_A_1_), .B(add_regs[29]), .CI(
        intadd_25_n5), .CO(intadd_25_n4), .S(intadd_25_SUM_1_) );
  ADFM1SA intadd_25_U6 ( .A(intadd_25_A_0_), .B(add_regs[28]), .CI(
        intadd_25_CI), .CO(intadd_25_n5), .S(intadd_25_SUM_0_) );
  DFQRM1SA shift_regs_reg_11__7_ ( .D(shift_regs[87]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[95]) );
  DFQRM1SA shift_regs_reg_11__6_ ( .D(shift_regs[86]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[94]) );
  DFQRM1SA shift_regs_reg_10__6_ ( .D(shift_regs[78]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[86]) );
  DFQRM1SA shift_regs_reg_10__5_ ( .D(shift_regs[77]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[85]) );
  DFQRM1SA shift_regs_reg_11__4_ ( .D(shift_regs[84]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[92]) );
  DFQRM1SA shift_regs_reg_10__4_ ( .D(shift_regs[76]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[84]) );
  DFQRM1SA shift_regs_reg_11__3_ ( .D(shift_regs[83]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[91]) );
  DFQRM1SA shift_regs_reg_10__3_ ( .D(shift_regs[75]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[83]) );
  DFQRM1SA shift_regs_reg_11__2_ ( .D(shift_regs[82]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[90]) );
  DFQRM1SA shift_regs_reg_10__2_ ( .D(shift_regs[74]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[82]) );
  DFQRM1SA shift_regs_reg_11__1_ ( .D(shift_regs[81]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[89]) );
  DFQRM1SA shift_regs_reg_10__1_ ( .D(shift_regs[73]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[81]) );
  DFQRM1SA shift_regs_reg_12__7_ ( .D(shift_regs[95]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[103]) );
  DFQRM1SA shift_regs_reg_9__7_ ( .D(shift_regs[71]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[79]) );
  DFQRM1SA shift_regs_reg_12__6_ ( .D(shift_regs[94]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[102]) );
  DFQRM1SA shift_regs_reg_9__6_ ( .D(shift_regs[70]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[78]) );
  DFQRM1SA shift_regs_reg_12__5_ ( .D(shift_regs[93]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[101]) );
  DFQRM1SA shift_regs_reg_9__5_ ( .D(shift_regs[69]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[77]) );
  DFQRM1SA shift_regs_reg_12__4_ ( .D(shift_regs[92]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[100]) );
  DFQRM1SA shift_regs_reg_9__4_ ( .D(shift_regs[68]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[76]) );
  DFQRM1SA shift_regs_reg_9__3_ ( .D(shift_regs[67]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[75]) );
  DFQRM1SA shift_regs_reg_12__2_ ( .D(shift_regs[90]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[98]) );
  DFQRM1SA shift_regs_reg_9__2_ ( .D(shift_regs[66]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[74]) );
  DFQRM1SA shift_regs_reg_12__1_ ( .D(shift_regs[89]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[97]) );
  DFQRM1SA shift_regs_reg_9__1_ ( .D(shift_regs[65]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[73]) );
  DFQRM1SA shift_regs_reg_12__0_ ( .D(shift_regs[88]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[96]) );
  DFQRM1SA shift_regs_reg_9__0_ ( .D(shift_regs[64]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[72]) );
  DFQRM1SA shift_regs_reg_13__7_ ( .D(shift_regs[103]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[111]) );
  DFQRM1SA shift_regs_reg_8__7_ ( .D(shift_regs[63]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[71]) );
  DFQRM1SA shift_regs_reg_13__6_ ( .D(shift_regs[102]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[110]) );
  DFQRM1SA shift_regs_reg_8__6_ ( .D(shift_regs[62]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[70]) );
  DFQRM1SA shift_regs_reg_13__5_ ( .D(shift_regs[101]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[109]) );
  DFQRM1SA shift_regs_reg_8__5_ ( .D(shift_regs[61]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[69]) );
  DFQRM1SA shift_regs_reg_13__3_ ( .D(shift_regs[99]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[107]) );
  DFQRM1SA shift_regs_reg_8__3_ ( .D(shift_regs[59]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[67]) );
  DFQRM1SA shift_regs_reg_13__2_ ( .D(shift_regs[98]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[106]) );
  DFQRM1SA shift_regs_reg_8__2_ ( .D(shift_regs[58]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[66]) );
  DFQRM1SA shift_regs_reg_8__1_ ( .D(shift_regs[57]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[65]) );
  DFQRM1SA shift_regs_reg_13__0_ ( .D(shift_regs[96]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[104]) );
  DFQRM1SA shift_regs_reg_8__0_ ( .D(shift_regs[56]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[64]) );
  DFQRM1SA shift_regs_reg_14__7_ ( .D(shift_regs[111]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[119]) );
  DFQRM1SA shift_regs_reg_7__7_ ( .D(shift_regs[55]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[63]) );
  DFQRM1SA shift_regs_reg_14__6_ ( .D(shift_regs[110]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[118]) );
  DFQRM1SA shift_regs_reg_7__6_ ( .D(shift_regs[54]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[62]) );
  DFQRM1SA shift_regs_reg_14__5_ ( .D(shift_regs[109]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[117]) );
  DFQRM1SA shift_regs_reg_7__5_ ( .D(shift_regs[53]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[61]) );
  DFQRM1SA shift_regs_reg_14__4_ ( .D(shift_regs[108]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[116]) );
  DFQRM1SA shift_regs_reg_7__4_ ( .D(shift_regs[52]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[60]) );
  DFQRM1SA shift_regs_reg_14__3_ ( .D(shift_regs[107]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[115]) );
  DFQRM1SA shift_regs_reg_7__3_ ( .D(shift_regs[51]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[59]) );
  DFQRM1SA shift_regs_reg_14__2_ ( .D(shift_regs[106]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[114]) );
  DFQRM1SA shift_regs_reg_7__2_ ( .D(shift_regs[50]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[58]) );
  DFQRM1SA shift_regs_reg_14__1_ ( .D(shift_regs[105]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[113]) );
  DFQRM1SA shift_regs_reg_7__1_ ( .D(shift_regs[49]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[57]) );
  DFQRM1SA shift_regs_reg_14__0_ ( .D(shift_regs[104]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[112]) );
  DFQRM1SA shift_regs_reg_7__0_ ( .D(shift_regs[48]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[56]) );
  DFQRM1SA shift_regs_reg_15__7_ ( .D(shift_regs[119]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[127]) );
  DFQRM1SA shift_regs_reg_6__7_ ( .D(shift_regs[47]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[55]) );
  DFQRM1SA shift_regs_reg_15__6_ ( .D(shift_regs[118]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[126]) );
  DFQRM1SA shift_regs_reg_6__6_ ( .D(shift_regs[46]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[54]) );
  DFQRM1SA shift_regs_reg_15__5_ ( .D(shift_regs[117]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[125]) );
  DFQRM1SA shift_regs_reg_6__5_ ( .D(shift_regs[45]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[53]) );
  DFQRM1SA shift_regs_reg_15__4_ ( .D(shift_regs[116]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[124]) );
  DFQRM1SA shift_regs_reg_6__4_ ( .D(shift_regs[44]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[52]) );
  DFQRM1SA shift_regs_reg_15__3_ ( .D(shift_regs[115]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[123]) );
  DFQRM1SA shift_regs_reg_6__3_ ( .D(shift_regs[43]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[51]) );
  DFQRM1SA shift_regs_reg_15__2_ ( .D(shift_regs[114]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[122]) );
  DFQRM1SA shift_regs_reg_6__2_ ( .D(shift_regs[42]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[50]) );
  DFQRM1SA shift_regs_reg_15__1_ ( .D(shift_regs[113]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[121]) );
  DFQRM1SA shift_regs_reg_6__1_ ( .D(shift_regs[41]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[49]) );
  DFQRM1SA shift_regs_reg_15__0_ ( .D(shift_regs[112]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[120]) );
  DFQRM1SA shift_regs_reg_16__7_ ( .D(shift_regs[127]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[135]) );
  DFQRM1SA shift_regs_reg_5__7_ ( .D(shift_regs[39]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[47]) );
  DFQRM1SA shift_regs_reg_16__6_ ( .D(shift_regs[126]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[134]) );
  DFQRM1SA shift_regs_reg_5__6_ ( .D(shift_regs[38]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[46]) );
  DFQRM1SA shift_regs_reg_16__5_ ( .D(shift_regs[125]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[133]) );
  DFQRM1SA shift_regs_reg_5__5_ ( .D(shift_regs[37]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[45]) );
  DFQRM1SA shift_regs_reg_16__4_ ( .D(shift_regs[124]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[132]) );
  DFQRM1SA shift_regs_reg_5__4_ ( .D(shift_regs[36]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[44]) );
  DFQRM1SA shift_regs_reg_16__3_ ( .D(shift_regs[123]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[131]) );
  DFQRM1SA shift_regs_reg_5__3_ ( .D(shift_regs[35]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[43]) );
  DFQRM1SA shift_regs_reg_16__2_ ( .D(shift_regs[122]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[130]) );
  DFQRM1SA shift_regs_reg_16__0_ ( .D(shift_regs[120]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[128]) );
  DFQRM1SA shift_regs_reg_5__0_ ( .D(shift_regs[32]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[40]) );
  DFQRM1SA shift_regs_reg_17__7_ ( .D(shift_regs[135]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[143]) );
  DFQRM1SA shift_regs_reg_4__7_ ( .D(shift_regs[31]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[39]) );
  DFQRM1SA shift_regs_reg_17__6_ ( .D(shift_regs[134]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[142]) );
  DFQRM1SA shift_regs_reg_4__6_ ( .D(shift_regs[30]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[38]) );
  DFQRM1SA shift_regs_reg_17__5_ ( .D(shift_regs[133]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[141]) );
  DFQRM1SA shift_regs_reg_4__5_ ( .D(shift_regs[29]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[37]) );
  DFQRM1SA shift_regs_reg_17__4_ ( .D(shift_regs[132]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[140]) );
  DFQRM1SA shift_regs_reg_17__3_ ( .D(shift_regs[131]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[139]) );
  DFQRM1SA shift_regs_reg_4__3_ ( .D(shift_regs[27]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[35]) );
  DFQRM1SA shift_regs_reg_17__2_ ( .D(shift_regs[130]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[138]) );
  DFQRM1SA shift_regs_reg_4__2_ ( .D(shift_regs[26]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[34]) );
  DFQRM1SA shift_regs_reg_17__1_ ( .D(shift_regs[129]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[137]) );
  DFQRM1SA shift_regs_reg_4__1_ ( .D(shift_regs[25]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[33]) );
  DFQRM1SA shift_regs_reg_17__0_ ( .D(shift_regs[128]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[136]) );
  DFQRM1SA shift_regs_reg_4__0_ ( .D(shift_regs[24]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[32]) );
  DFQRM1SA shift_regs_reg_18__7_ ( .D(shift_regs[143]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[151]) );
  DFQRM1SA shift_regs_reg_3__7_ ( .D(shift_regs[23]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[31]) );
  DFQRM1SA shift_regs_reg_18__5_ ( .D(shift_regs[141]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[149]) );
  DFQRM1SA shift_regs_reg_3__5_ ( .D(shift_regs[21]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[29]) );
  DFQRM1SA shift_regs_reg_18__3_ ( .D(shift_regs[139]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[147]) );
  DFQRM1SA shift_regs_reg_3__3_ ( .D(shift_regs[19]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[27]) );
  DFQRM1SA shift_regs_reg_18__2_ ( .D(shift_regs[138]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[146]) );
  DFQRM1SA shift_regs_reg_3__2_ ( .D(shift_regs[18]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[26]) );
  DFQRM1SA shift_regs_reg_18__1_ ( .D(shift_regs[137]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[145]) );
  DFQRM1SA shift_regs_reg_3__1_ ( .D(shift_regs[17]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[25]) );
  DFQRM1SA shift_regs_reg_18__0_ ( .D(shift_regs[136]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[144]) );
  DFQRM1SA shift_regs_reg_3__0_ ( .D(shift_regs[16]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[24]) );
  DFQRM1SA shift_regs_reg_19__7_ ( .D(shift_regs[151]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[159]) );
  DFQRM1SA shift_regs_reg_2__7_ ( .D(shift_regs[15]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[23]) );
  DFQRM1SA shift_regs_reg_19__6_ ( .D(shift_regs[150]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[158]) );
  DFQRM1SA shift_regs_reg_2__6_ ( .D(shift_regs[14]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[22]) );
  DFQRM1SA shift_regs_reg_19__5_ ( .D(shift_regs[149]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[157]) );
  DFQRM1SA shift_regs_reg_2__5_ ( .D(shift_regs[13]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[21]) );
  DFQRM1SA shift_regs_reg_2__4_ ( .D(shift_regs[12]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[20]) );
  DFQRM1SA shift_regs_reg_19__2_ ( .D(shift_regs[146]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[154]) );
  DFQRM1SA shift_regs_reg_2__2_ ( .D(shift_regs[10]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[18]) );
  DFQRM1SA shift_regs_reg_19__1_ ( .D(shift_regs[145]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[153]) );
  DFQRM1SA shift_regs_reg_2__1_ ( .D(shift_regs[9]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[17]) );
  DFQRM1SA shift_regs_reg_19__0_ ( .D(shift_regs[144]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[152]) );
  DFQRM1SA shift_regs_reg_2__0_ ( .D(shift_regs[8]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[16]) );
  DFQRM1SA shift_regs_reg_20__7_ ( .D(shift_regs[159]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[167]) );
  DFQRM1SA shift_regs_reg_1__7_ ( .D(shift_regs[7]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[15]) );
  DFQRM1SA shift_regs_reg_20__6_ ( .D(shift_regs[158]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[166]) );
  DFQRM1SA shift_regs_reg_1__6_ ( .D(shift_regs[6]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[14]) );
  DFQRM1SA shift_regs_reg_20__5_ ( .D(shift_regs[157]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[165]) );
  DFQRM1SA shift_regs_reg_1__5_ ( .D(shift_regs[5]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[13]) );
  DFQRM1SA shift_regs_reg_20__4_ ( .D(shift_regs[156]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[164]) );
  DFQRM1SA shift_regs_reg_1__4_ ( .D(shift_regs[4]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[12]) );
  DFQRM1SA shift_regs_reg_20__3_ ( .D(shift_regs[155]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[163]) );
  DFQRM1SA shift_regs_reg_1__3_ ( .D(shift_regs[3]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[11]) );
  DFQRM1SA shift_regs_reg_1__2_ ( .D(shift_regs[2]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[10]) );
  DFQRM1SA shift_regs_reg_20__0_ ( .D(shift_regs[152]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[160]) );
  DFQRM1SA shift_regs_reg_1__0_ ( .D(shift_regs[0]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[8]) );
  DFQRM1SA shift_regs_reg_21__7_ ( .D(shift_regs[167]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[175]) );
  DFQRM1SA shift_regs_reg_0__7_ ( .D(input_data[7]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[7]) );
  DFQRM1SA shift_regs_reg_21__6_ ( .D(shift_regs[166]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[174]) );
  DFQRM1SA shift_regs_reg_0__6_ ( .D(input_data[6]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[6]) );
  DFQRM1SA shift_regs_reg_21__5_ ( .D(shift_regs[165]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[173]) );
  DFQRM1SA shift_regs_reg_0__5_ ( .D(input_data[5]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[5]) );
  DFQRM1SA shift_regs_reg_21__4_ ( .D(shift_regs[164]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[172]) );
  DFQRM1SA shift_regs_reg_0__4_ ( .D(input_data[4]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[4]) );
  DFQRM1SA shift_regs_reg_21__3_ ( .D(shift_regs[163]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[171]) );
  DFQRM1SA shift_regs_reg_0__3_ ( .D(input_data[3]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[3]) );
  DFQRM1SA shift_regs_reg_21__2_ ( .D(shift_regs[162]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[170]) );
  DFQRM1SA shift_regs_reg_0__2_ ( .D(input_data[2]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[2]) );
  DFQRM1SA shift_regs_reg_21__1_ ( .D(shift_regs[161]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[169]) );
  DFQRM1SA shift_regs_reg_0__1_ ( .D(input_data[1]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[1]) );
  DFQRM1SA shift_regs_reg_0__0_ ( .D(input_data[0]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[0]) );
  ADFM1SA intadd_2_U8 ( .A(add_regs[73]), .B(intadd_2_B_1_), .CI(intadd_2_n8), 
        .CO(intadd_2_n7), .S(intadd_2_SUM_1_) );
  ADFM1SA intadd_3_U8 ( .A(add_regs[68]), .B(intadd_3_B_0_), .CI(intadd_3_CI), 
        .CO(intadd_3_n7), .S(intadd_3_SUM_0_) );
  ADFM1SA intadd_32_U3 ( .A(intadd_32_A_2_), .B(intadd_32_B_2_), .CI(
        intadd_32_n3), .CO(intadd_32_n2), .S(intadd_32_SUM_2_) );
  DFQRM1SA shift_regs_reg_11__0_ ( .D(shift_regs[80]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[88]) );
  DFQRM1SA shift_regs_reg_10__0_ ( .D(shift_regs[72]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[80]) );
  DFQRM1SA shift_regs_reg_13__4_ ( .D(shift_regs[100]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[108]) );
  DFQRM1SA shift_regs_reg_8__4_ ( .D(shift_regs[60]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[68]) );
  DFQRM1SA shift_regs_reg_16__1_ ( .D(shift_regs[121]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[129]) );
  DFQRM1SA shift_regs_reg_5__1_ ( .D(shift_regs[33]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[41]) );
  DFQRM1SA shift_regs_reg_18__4_ ( .D(shift_regs[140]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[148]) );
  DFQRM1SA shift_regs_reg_3__4_ ( .D(shift_regs[20]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[28]) );
  DFQRM1SA shift_regs_reg_19__3_ ( .D(shift_regs[147]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[155]) );
  DFQRM1SA shift_regs_reg_2__3_ ( .D(shift_regs[11]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[19]) );
  DFQRM1SA shift_regs_reg_20__1_ ( .D(shift_regs[153]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[161]) );
  DFQRM1SA shift_regs_reg_1__1_ ( .D(shift_regs[1]), .CK(CLK_Filter), .RB(
        rst_n), .Q(shift_regs[9]) );
  ADFM1SA intadd_26_U3 ( .A(intadd_26_A_2_), .B(intadd_26_B_2_), .CI(
        intadd_26_n3), .CO(intadd_26_n2), .S(intadd_26_SUM_2_) );
  ADFM1SA intadd_27_U3 ( .A(intadd_27_A_2_), .B(intadd_27_B_2_), .CI(
        intadd_27_n3), .CO(intadd_27_n2), .S(intadd_27_SUM_2_) );
  ADFM1SA intadd_17_U3 ( .A(intadd_17_A_3_), .B(intadd_17_B_3_), .CI(
        intadd_17_n3), .CO(intadd_17_n2), .S(intadd_17_SUM_3_) );
  ADFM1SA intadd_34_U2 ( .A(intadd_27_SUM_1_), .B(intadd_34_B_2_), .CI(
        intadd_34_n2), .CO(intadd_34_n1), .S(intadd_18_A_4_) );
  ADFM1SA intadd_18_U3 ( .A(intadd_18_A_3_), .B(intadd_18_B_3_), .CI(
        intadd_18_n3), .CO(intadd_18_n2), .S(intadd_18_SUM_3_) );
  ADFM1SA intadd_19_U3 ( .A(intadd_19_A_3_), .B(intadd_33_n1), .CI(
        intadd_19_n3), .CO(intadd_19_n2), .S(intadd_19_SUM_3_) );
  ADFM1SA intadd_17_U4 ( .A(intadd_17_A_2_), .B(intadd_17_B_2_), .CI(
        intadd_17_n4), .CO(intadd_17_n3), .S(intadd_17_SUM_2_) );
  ADFM1SA intadd_20_U3 ( .A(intadd_20_A_3_), .B(intadd_18_SUM_1_), .CI(
        intadd_20_n3), .CO(intadd_20_n2), .S(intadd_20_SUM_3_) );
  ADFM1SA intadd_18_U4 ( .A(intadd_17_SUM_1_), .B(intadd_18_B_2_), .CI(
        intadd_18_n4), .CO(intadd_18_n3), .S(intadd_18_SUM_2_) );
  ADFM1SA intadd_21_U3 ( .A(intadd_21_A_3_), .B(intadd_19_SUM_1_), .CI(
        intadd_21_n3), .CO(intadd_21_n2), .S(intadd_21_SUM_3_) );
  ADFM1SA intadd_19_U4 ( .A(intadd_19_A_2_), .B(intadd_19_B_2_), .CI(
        intadd_19_n4), .CO(intadd_19_n3), .S(intadd_19_SUM_2_) );
  ADFM1SA intadd_22_U3 ( .A(intadd_22_A_3_), .B(intadd_20_SUM_1_), .CI(
        intadd_22_n3), .CO(intadd_22_n2), .S(intadd_22_SUM_3_) );
  ADFM1SA intadd_20_U4 ( .A(intadd_20_A_2_), .B(intadd_20_B_2_), .CI(
        intadd_20_n4), .CO(intadd_20_n3), .S(intadd_20_SUM_2_) );
  ADFM1SA intadd_23_U3 ( .A(intadd_23_A_3_), .B(intadd_21_SUM_1_), .CI(
        intadd_23_n3), .CO(intadd_23_n2), .S(intadd_23_SUM_3_) );
  ADFM1SA intadd_21_U4 ( .A(intadd_21_A_2_), .B(intadd_21_B_2_), .CI(
        intadd_21_n4), .CO(intadd_21_n3), .S(intadd_21_SUM_2_) );
  ADFM1SA intadd_24_U3 ( .A(intadd_24_A_3_), .B(intadd_22_SUM_1_), .CI(
        intadd_24_n3), .CO(intadd_24_n2), .S(intadd_24_SUM_3_) );
  ADFM1SA intadd_22_U4 ( .A(intadd_20_SUM_0_), .B(intadd_22_B_2_), .CI(
        intadd_22_n4), .CO(intadd_22_n3), .S(intadd_22_SUM_2_) );
  ADFM1SA intadd_28_U3 ( .A(intadd_28_A_2_), .B(intadd_23_SUM_1_), .CI(
        intadd_28_n3), .CO(intadd_28_n2), .S(intadd_28_SUM_2_) );
  ADFM1SA intadd_23_U4 ( .A(intadd_21_SUM_0_), .B(intadd_23_B_2_), .CI(
        intadd_23_n4), .CO(intadd_23_n3), .S(intadd_23_SUM_2_) );
  ADFM1SA intadd_29_U3 ( .A(intadd_24_SUM_1_), .B(intadd_23_SUM_0_), .CI(
        intadd_29_n3), .CO(intadd_29_n2), .S(intadd_29_SUM_2_) );
  ADFM1SA intadd_24_U4 ( .A(intadd_24_A_2_), .B(intadd_22_SUM_0_), .CI(
        intadd_24_n4), .CO(intadd_24_n3), .S(intadd_24_SUM_2_) );
  ADFM1SA intadd_28_U4 ( .A(intadd_28_A_1_), .B(intadd_28_B_1_), .CI(
        intadd_28_n4), .CO(intadd_28_n3), .S(intadd_28_SUM_1_) );
  ADFM1SA intadd_29_U4 ( .A(intadd_29_A_1_), .B(intadd_29_B_1_), .CI(
        intadd_29_n4), .CO(intadd_29_n3), .S(intadd_29_SUM_1_) );
  ADFM1SA intadd_28_U5 ( .A(order[58]), .B(order[88]), .CI(order[31]), .CO(
        intadd_28_n4), .S(intadd_28_SUM_0_) );
  ADFM1SA intadd_24_U6 ( .A(order[11]), .B(order[119]), .CI(order[2]), .CO(
        intadd_24_n5), .S(intadd_24_SUM_0_) );
  ADFM1SA intadd_29_U5 ( .A(order[44]), .B(order[71]), .CI(order[103]), .CO(
        intadd_29_n4), .S(intadd_29_SUM_0_) );
  DFQRM1SA order_reg_1__1_ ( .D(N101), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[9]) );
  DFQRM1SA order_reg_0__1_ ( .D(add_regs[0]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[0]) );
  DFQRM1SA order_reg_9__1_ ( .D(N206), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[117]) );
  DFQRM1SA order_reg_6__1_ ( .D(N158), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[70]) );
  ADFM1SA intadd_26_U4 ( .A(intadd_26_A_1_), .B(intadd_26_B_1_), .CI(
        intadd_26_n4), .CO(intadd_26_n3), .S(intadd_26_SUM_1_) );
  ADFM1SA intadd_27_U4 ( .A(intadd_27_A_1_), .B(intadd_27_B_1_), .CI(
        intadd_27_n4), .CO(intadd_27_n3), .S(intadd_27_SUM_1_) );
  ADFM1SA intadd_34_U3 ( .A(intadd_34_A_1_), .B(intadd_34_B_1_), .CI(
        intadd_34_n3), .CO(intadd_34_n2), .S(intadd_17_A_2_) );
  ADFM1SA intadd_33_U2 ( .A(intadd_33_A_2_), .B(intadd_17_SUM_0_), .CI(
        intadd_33_n2), .CO(intadd_33_n1), .S(intadd_20_A_3_) );
  ADFM1SA intadd_17_U5 ( .A(intadd_17_A_1_), .B(intadd_17_B_1_), .CI(
        intadd_17_n5), .CO(intadd_17_n4), .S(intadd_17_SUM_1_) );
  ADFM1SA intadd_18_U5 ( .A(intadd_18_A_1_), .B(intadd_18_B_1_), .CI(
        intadd_18_n5), .CO(intadd_18_n4), .S(intadd_18_SUM_1_) );
  ADFM1SA intadd_19_U5 ( .A(intadd_19_A_1_), .B(intadd_19_B_1_), .CI(
        intadd_19_n5), .CO(intadd_19_n4), .S(intadd_19_SUM_1_) );
  ADFM1SA intadd_20_U5 ( .A(intadd_20_A_1_), .B(intadd_20_B_1_), .CI(
        intadd_20_n5), .CO(intadd_20_n4), .S(intadd_20_SUM_1_) );
  ADFM1SA intadd_33_U3 ( .A(order[94]), .B(order[64]), .CI(intadd_33_n3), .CO(
        intadd_33_n2), .S(intadd_20_A_2_) );
  ADFM1SA intadd_21_U5 ( .A(intadd_21_A_1_), .B(intadd_21_B_1_), .CI(
        intadd_21_n5), .CO(intadd_21_n4), .S(intadd_21_SUM_1_) );
  ADFM1SA intadd_22_U5 ( .A(order[61]), .B(intadd_22_B_1_), .CI(intadd_22_n5), 
        .CO(intadd_22_n4), .S(intadd_22_SUM_1_) );
  ADFM1SA intadd_20_U6 ( .A(order[49]), .B(order[123]), .CI(order[76]), .CO(
        intadd_20_n5), .S(intadd_20_SUM_0_) );
  ADFM1SA intadd_23_U5 ( .A(order[60]), .B(order[33]), .CI(intadd_23_n5), .CO(
        intadd_23_n4), .S(intadd_23_SUM_1_) );
  ADFM1SA intadd_21_U6 ( .A(order[48]), .B(order[75]), .CI(order[107]), .CO(
        intadd_21_n5), .S(intadd_21_SUM_0_) );
  ADFM1SA intadd_24_U5 ( .A(order[59]), .B(intadd_24_B_1_), .CI(intadd_24_n5), 
        .CO(intadd_24_n4), .S(intadd_24_SUM_1_) );
  ADFM1SA intadd_23_U6 ( .A(order[46]), .B(order[73]), .CI(order[105]), .CO(
        intadd_23_n5), .S(intadd_23_SUM_0_) );
  ADFM1SA intadd_22_U6 ( .A(order[22]), .B(order[121]), .CI(order[47]), .CO(
        intadd_22_n5), .S(intadd_22_SUM_0_) );
  DFQRM1SA order_reg_9__2_ ( .D(N207), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[118]) );
  DFQRM1SA order_reg_5__2_ ( .D(N144), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[57]) );
  DFQRM1SA order_reg_3__2_ ( .D(N115), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[30]) );
  DFQRM1SA order_reg_1__2_ ( .D(N102), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[10]) );
  DFQRM1SA order_reg_0__2_ ( .D(add_regs[1]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[1]) );
  ADFM1SA intadd_26_U5 ( .A(order[55]), .B(order[41]), .CI(order[82]), .CO(
        intadd_26_n4), .S(intadd_26_SUM_0_) );
  DFQRM1SA order_reg_10__14_ ( .D(add_regs[87]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[139]) );
  DFQRM1SA order_reg_10__13_ ( .D(add_regs[86]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[138]) );
  ADFM1SA intadd_27_U5 ( .A(order[54]), .B(order[128]), .CI(order[81]), .CO(
        intadd_27_n4), .S(intadd_27_SUM_0_) );
  ADFM1SA intadd_34_U4 ( .A(order[39]), .B(order[28]), .CI(order[19]), .CO(
        intadd_34_n3), .S(intadd_34_SUM_0_) );
  DFQRM1SA order_reg_10__12_ ( .D(add_regs[85]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[137]) );
  ADFM1SA intadd_17_U6 ( .A(order[38]), .B(order[27]), .CI(order[18]), .CO(
        intadd_17_n5), .S(intadd_17_SUM_0_) );
  DFQRM1SA order_reg_10__11_ ( .D(add_regs[84]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[136]) );
  ADFM1SA intadd_18_U6 ( .A(order[26]), .B(order[125]), .CI(order[51]), .CO(
        intadd_18_n5), .S(intadd_18_SUM_0_) );
  DFQRM1SA order_reg_10__10_ ( .D(add_regs[83]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[135]) );
  ADFM1SA intadd_19_U6 ( .A(order[16]), .B(order[93]), .CI(order[7]), .CO(
        intadd_19_n5), .S(intadd_19_SUM_0_) );
  ADFM1SA intadd_33_U4 ( .A(order[77]), .B(order[109]), .CI(order[133]), .CO(
        intadd_33_n3), .S(intadd_33_SUM_0_) );
  DFQRM1SA order_reg_10__7_ ( .D(add_regs[80]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[132]) );
  DFQRM1SA order_reg_2__5_ ( .D(add_regs[17]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[22]) );
  DFQRM1SA order_reg_0__5_ ( .D(add_regs[4]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[4]) );
  DFQRM1SA order_reg_0__4_ ( .D(add_regs[3]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[3]) );
  DFQRM1SA order_reg_2__4_ ( .D(add_regs[16]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[21]) );
  DFQRM1SA order_reg_2__12_ ( .D(add_regs[24]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[29]) );
  DFQRM1SA order_reg_2__11_ ( .D(add_regs[23]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[28]) );
  DFQRM1SA order_reg_2__10_ ( .D(add_regs[22]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[27]) );
  DFQRM1SA order_reg_2__9_ ( .D(add_regs[21]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[26]) );
  DFQRM1SA order_reg_0__9_ ( .D(add_regs[8]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[8]) );
  DFQRM1SA order_reg_10__9_ ( .D(add_regs[82]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[134]) );
  DFQRM1SA order_reg_0__8_ ( .D(add_regs[7]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[7]) );
  DFQRM1SA order_reg_2__8_ ( .D(add_regs[20]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[25]) );
  DFQRM1SA order_reg_0__7_ ( .D(add_regs[6]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[6]) );
  DFQRM1SA order_reg_2__7_ ( .D(add_regs[19]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[24]) );
  DFQRM1SA order_reg_10__8_ ( .D(add_regs[81]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[133]) );
  DFQRM1SA order_reg_0__6_ ( .D(add_regs[5]), .CK(CLK_Filter), .RB(rst_n), .Q(
        order[5]) );
  DFQRM1SA order_reg_2__6_ ( .D(add_regs[18]), .CK(CLK_Filter), .RB(rst_n), 
        .Q(order[23]) );
  INVM1S U6 ( .A(1'b1), .Z(output_data[19]) );
  ADFM1SA U8 ( .A(order[5]), .B(order[122]), .CI(order[23]), .CO(n53), .S(n51)
         );
  ADFM1SA U9 ( .A(order[34]), .B(order[91]), .CI(order[14]), .CO(
        intadd_21_B_1_), .S(n49) );
  ADFM1SA U10 ( .A(order[6]), .B(order[92]), .CI(order[24]), .CO(
        intadd_20_A_1_), .S(n54) );
  ADFM1SA U11 ( .A(order[35]), .B(order[62]), .CI(order[15]), .CO(
        intadd_20_B_1_), .S(n52) );
  ADFM1SA U12 ( .A(order[25]), .B(order[124]), .CI(order[50]), .CO(
        intadd_19_B_1_), .S(n55) );
  ADFM1SA U13 ( .A(order[78]), .B(order[110]), .CI(order[134]), .CO(n58), .S(
        n57) );
  ADFM1SA U14 ( .A(order[37]), .B(order[8]), .CI(order[17]), .CO(
        intadd_18_B_1_), .S(intadd_19_A_1_) );
  ADFM1SA U15 ( .A(order[52]), .B(order[126]), .CI(order[79]), .CO(
        intadd_17_B_1_), .S(intadd_33_A_2_) );
  ADFM1SA U16 ( .A(order[53]), .B(order[127]), .CI(order[80]), .CO(
        intadd_34_B_1_), .S(n60) );
  ADFM1SA U17 ( .A(order[96]), .B(order[66]), .CI(n138), .CO(n61), .S(n59) );
  ADFM1SA U18 ( .A(order[40]), .B(order[29]), .CI(order[20]), .CO(
        intadd_27_A_1_), .S(n62) );
  ADFM1SA U19 ( .A(order[68]), .B(order[98]), .CI(order[114]), .CO(
        intadd_26_B_1_), .S(n65) );
  ADFM1SA U20 ( .A(order[32]), .B(order[89]), .CI(order[12]), .CO(n47), .S(
        intadd_28_B_1_) );
  ADFM1SA U21 ( .A(order[3]), .B(order[120]), .CI(order[21]), .CO(n46), .S(
        intadd_28_A_1_) );
  ADFM1SA U22 ( .A(order[13]), .B(order[90]), .CI(order[4]), .CO(n50), .S(
        intadd_24_A_2_) );
  ADFM1SA U23 ( .A(n48), .B(n47), .CI(n46), .CO(intadd_23_B_2_), .S(
        intadd_28_A_2_) );
  ADFM1SA U24 ( .A(n51), .B(n50), .CI(n49), .CO(intadd_22_B_2_), .S(
        intadd_24_A_3_) );
  ADFM1SA U25 ( .A(order[63]), .B(order[36]), .CI(n139), .CO(n56), .S(
        intadd_21_A_2_) );
  ADFM1SA U26 ( .A(n54), .B(n53), .CI(n52), .CO(intadd_21_B_2_), .S(
        intadd_23_A_3_) );
  ADFM1SA U27 ( .A(n55), .B(intadd_33_SUM_0_), .CI(intadd_19_SUM_0_), .CO(
        intadd_20_B_2_), .S(intadd_22_A_3_) );
  ADFM1SA U28 ( .A(n57), .B(n56), .CI(intadd_18_SUM_0_), .CO(intadd_19_B_2_), 
        .S(intadd_21_A_3_) );
  ADFM1SA U29 ( .A(order[95]), .B(order[65]), .CI(n58), .CO(intadd_18_B_2_), 
        .S(intadd_19_A_2_) );
  ADFM1SA U30 ( .A(n60), .B(n59), .CI(intadd_34_SUM_0_), .CO(intadd_18_B_3_), 
        .S(intadd_19_A_3_) );
  ADFM1SA U31 ( .A(order[97]), .B(order[67]), .CI(n137), .CO(intadd_34_B_2_), 
        .S(intadd_17_B_2_) );
  ADFM1SA U32 ( .A(n62), .B(n61), .CI(intadd_27_SUM_0_), .CO(intadd_17_B_3_), 
        .S(intadd_18_A_3_) );
  ADFM1SA U33 ( .A(n65), .B(n64), .CI(intadd_26_SUM_0_), .CO(n63), .S(
        intadd_17_A_3_) );
  ADFM1SA U34 ( .A(order[83]), .B(order[99]), .CI(order[115]), .CO(n67), .S(
        intadd_27_B_2_) );
  ADFM1SA U35 ( .A(order[69]), .B(order[56]), .CI(n69), .CO(n66), .S(
        intadd_27_A_2_) );
  ADFM1SA U36 ( .A(add_regs[36]), .B(add_regs[38]), .CI(add_regs[34]), .CO(n30), .S(n80) );
  ADFM1SA U37 ( .A(add_regs[54]), .B(n98), .CI(intadd_32_B_0_), .CO(
        intadd_32_B_3_), .S(intadd_32_A_2_) );
  ADFM1SA U38 ( .A(add_regs[67]), .B(add_regs[71]), .CI(n128), .CO(
        intadd_3_A_3_), .S(intadd_3_B_2_) );
  ADFM1SA U39 ( .A(add_regs[72]), .B(n127), .CI(add_regs[68]), .CO(
        intadd_3_B_4_), .S(intadd_3_B_3_) );
  ADFM1SA U40 ( .A(N207), .B(add_regs[78]), .CI(intadd_2_B_2_), .CO(n154), .S(
        n155) );
  ADFM1SA U41 ( .A(add_regs[73]), .B(add_regs[79]), .CI(n157), .CO(n152), .S(
        n153) );
  ADFM1SA U42 ( .A(order[30]), .B(order[10]), .CI(order[1]), .CO(
        intadd_29_A_1_), .S(n42) );
  ADFM1SA U43 ( .A(order[87]), .B(order[118]), .CI(order[57]), .CO(
        intadd_29_B_1_), .S(intadd_35_A_1_) );
  ADFM1SA U44 ( .A(order[45]), .B(order[72]), .CI(order[104]), .CO(
        intadd_24_B_1_), .S(n45) );
  ADFM1SA U45 ( .A(intadd_27_SUM_2_), .B(n63), .CI(intadd_26_SUM_1_), .CO(
        intadd_27_B_3_), .S(intadd_17_A_4_) );
  ADFM1SA U46 ( .A(order[84]), .B(order[100]), .CI(n136), .CO(n135), .S(
        intadd_26_B_2_) );
  ADFM1SA U47 ( .A(order[116]), .B(order[131]), .CI(order[140]), .CO(n134), 
        .S(n68) );
  ADFM1SA U48 ( .A(n68), .B(n67), .CI(n66), .CO(intadd_26_B_3_), .S(
        intadd_26_A_2_) );
  ADFM1SA U49 ( .A(add_regs[36]), .B(add_regs[37]), .CI(n27), .CO(
        intadd_1_B_3_), .S(intadd_1_A_2_) );
  ADFM1SA U50 ( .A(add_regs[38]), .B(n29), .CI(n90), .CO(intadd_1_B_4_), .S(
        intadd_1_A_3_) );
  ADFM1SA U51 ( .A(n86), .B(n85), .CI(n84), .CO(n83), .S(n87) );
  ADFM1SA U52 ( .A(add_regs[40]), .B(n31), .CI(n30), .CO(intadd_1_B_6_), .S(
        intadd_1_A_5_) );
  ADFM1SA U53 ( .A(n78), .B(n77), .CI(n76), .CO(n75), .S(n79) );
  ADFM1SA U54 ( .A(add_regs[56]), .B(n98), .CI(n100), .CO(n97), .S(n99) );
  ADFM1SA U55 ( .A(add_regs[63]), .B(n115), .CI(n114), .CO(n112), .S(n113) );
  ADFM1SA U56 ( .A(add_regs[64]), .B(n114), .CI(n110), .CO(n109), .S(n111) );
  ADFM1SA U57 ( .A(order[117]), .B(order[86]), .CI(n43), .CO(n41), .S(
        intadd_0_A_1_) );
  ADFM1SA U58 ( .A(n42), .B(n41), .CI(intadd_29_SUM_0_), .CO(intadd_35_B_2_), 
        .S(intadd_0_A_2_) );
  ADFM1SA U59 ( .A(intadd_28_SUM_0_), .B(n45), .CI(intadd_24_SUM_0_), .CO(n44), 
        .S(intadd_0_B_3_) );
  ADFM1SA U60 ( .A(intadd_29_SUM_2_), .B(n44), .CI(intadd_28_SUM_1_), .CO(
        intadd_0_B_5_), .S(intadd_0_A_4_) );
  MAOI22M1SA U61 ( .A1(n71), .A2(n72), .B1(n71), .B2(n72), .Z(intadd_1_A_7_)
         );
  MAOI22M1SA U62 ( .A1(add_regs[31]), .A2(n24), .B1(add_regs[31]), .B2(n24), 
        .Z(N125) );
  OA21M1SA U63 ( .A1(n35), .A2(n98), .B(intadd_32_CI), .Z(N161) );
  MAOI22M1SA U64 ( .A1(n118), .A2(n108), .B1(n118), .B2(n108), .Z(N177) );
  MAOI22M1SA U65 ( .A1(N189), .A2(n16), .B1(N189), .B2(n16), .Z(N193) );
  INVM1S U66 ( .A(intadd_25_n1), .Z(n23) );
  NR2M2S U67 ( .A(add_regs[30]), .B(n23), .Z(n24) );
  INVM1S U68 ( .A(add_regs[33]), .Z(n89) );
  NR2M1S U69 ( .A(N127), .B(n89), .Z(n26) );
  MAOI22M1SA U70 ( .A1(n26), .A2(add_regs[34]), .B1(n26), .B2(add_regs[34]), 
        .Z(N129) );
  INVM1S U71 ( .A(add_regs[35]), .Z(n88) );
  ND2M1S U72 ( .A(n88), .B(n89), .Z(n82) );
  NR2M1S U73 ( .A(n88), .B(n89), .Z(n81) );
  NR2B1M2S U74 ( .NA(n82), .B(n81), .Z(n28) );
  MAOI22M1SA U75 ( .A1(add_regs[36]), .A2(n28), .B1(add_regs[36]), .B2(n28), 
        .Z(intadd_1_A_1_) );
  INVM1S U76 ( .A(add_regs[42]), .Z(intadd_30_B_1_) );
  INVM1S U77 ( .A(add_regs[44]), .Z(intadd_30_B_3_) );
  NR2M1S U78 ( .A(N144), .B(add_regs[41]), .Z(n146) );
  ND2M1S U79 ( .A(n146), .B(intadd_30_B_1_), .Z(n145) );
  NR2M2S U80 ( .A(add_regs[43]), .B(n145), .Z(n144) );
  MAOI22M1SA U81 ( .A1(N144), .A2(intadd_30_B_3_), .B1(intadd_30_B_3_), .B2(
        N144), .Z(n10) );
  MAOI22M1SA U82 ( .A1(n144), .A2(n10), .B1(n144), .B2(n10), .Z(N148) );
  INVM1S U83 ( .A(add_regs[45]), .Z(n148) );
  ND2M1S U84 ( .A(intadd_30_n1), .B(n148), .Z(n147) );
  NR2M2S U85 ( .A(add_regs[46]), .B(n147), .Z(n32) );
  MAOI22M1SA U86 ( .A1(add_regs[47]), .A2(n32), .B1(add_regs[47]), .B2(n32), 
        .Z(N155) );
  INVM1S U87 ( .A(N158), .Z(intadd_32_A_1_) );
  INVM1S U88 ( .A(add_regs[49]), .Z(intadd_32_B_0_) );
  ND2M1S U89 ( .A(intadd_32_A_1_), .B(intadd_32_B_0_), .Z(n34) );
  MAOI22M1SA U90 ( .A1(add_regs[50]), .A2(n34), .B1(add_regs[50]), .B2(n34), 
        .Z(N160) );
  INVM1S U91 ( .A(add_regs[55]), .Z(intadd_31_CI) );
  INVM1S U92 ( .A(add_regs[56]), .Z(n104) );
  INVM1S U93 ( .A(add_regs[54]), .Z(n101) );
  AOI22M1S U94 ( .A1(add_regs[56]), .A2(add_regs[54]), .B1(n104), .B2(n101), 
        .Z(n12) );
  INVM1S U95 ( .A(add_regs[53]), .Z(n100) );
  ND2M1S U96 ( .A(intadd_31_CI), .B(n100), .Z(n95) );
  ND2M1S U97 ( .A(intadd_31_n1), .B(n95), .Z(n102) );
  OAI21M1S U98 ( .A1(intadd_31_n1), .A2(n95), .B(n102), .Z(n11) );
  MAOI22M1SA U99 ( .A1(n12), .A2(n11), .B1(n12), .B2(n11), .Z(N169) );
  NR2M1S U100 ( .A(N173), .B(add_regs[57]), .Z(n120) );
  INVM1S U101 ( .A(add_regs[58]), .Z(n114) );
  ND2M1S U102 ( .A(n120), .B(n114), .Z(n119) );
  NR2M1S U103 ( .A(add_regs[59]), .B(n119), .Z(n118) );
  INVM1S U104 ( .A(add_regs[60]), .Z(n108) );
  INVM1S U105 ( .A(add_regs[25]), .Z(intadd_25_A_0_) );
  INVM1S U106 ( .A(add_regs[27]), .Z(intadd_25_B_2_) );
  INVM1S U107 ( .A(N115), .Z(n70) );
  ND2M1S U108 ( .A(n70), .B(intadd_25_A_0_), .Z(n143) );
  NR2M2S U109 ( .A(add_regs[26]), .B(n143), .Z(n142) );
  AOI22M1S U110 ( .A1(N115), .A2(intadd_25_B_2_), .B1(add_regs[27]), .B2(n70), 
        .Z(n13) );
  MAOI22M1SA U111 ( .A1(n142), .A2(n13), .B1(n142), .B2(n13), .Z(N118) );
  INVM1S U112 ( .A(add_regs[62]), .Z(n106) );
  INVM1S U113 ( .A(add_regs[64]), .Z(n121) );
  OAI21M1S U114 ( .A1(n106), .A2(add_regs[63]), .B(n121), .Z(n14) );
  OAI31M1S U115 ( .A1(n106), .A2(add_regs[63]), .A3(n121), .B(n14), .Z(n15) );
  MAOI22M1SA U116 ( .A1(intadd_4_n1), .A2(n15), .B1(intadd_4_n1), .B2(n15), 
        .Z(N186) );
  INVM1S U117 ( .A(add_regs[63]), .Z(n123) );
  ND2M1S U118 ( .A(n106), .B(n123), .Z(n105) );
  ND2M1S U119 ( .A(intadd_4_n1), .B(n105), .Z(n122) );
  AO33M1SA U120 ( .A1(add_regs[63]), .A2(n121), .A3(intadd_4_n1), .B1(n123), 
        .B2(add_regs[64]), .B3(n122), .Z(N187) );
  NR2M1S U121 ( .A(N189), .B(add_regs[65]), .Z(n131) );
  INVM1S U122 ( .A(add_regs[66]), .Z(n125) );
  ND2M1S U123 ( .A(n131), .B(n125), .Z(n130) );
  NR2M2S U124 ( .A(add_regs[67]), .B(n130), .Z(n129) );
  INVM1S U125 ( .A(add_regs[68]), .Z(n39) );
  MAOI22M1SA U126 ( .A1(n129), .A2(n39), .B1(n129), .B2(n39), .Z(n16) );
  INVM1S U127 ( .A(add_regs[69]), .Z(n126) );
  INVM1S U128 ( .A(add_regs[72]), .Z(n132) );
  AOI22M1S U129 ( .A1(add_regs[72]), .A2(n126), .B1(add_regs[69]), .B2(n132), 
        .Z(n19) );
  INVM1S U130 ( .A(intadd_3_n1), .Z(n17) );
  ND2M1S U131 ( .A(add_regs[71]), .B(n39), .Z(n38) );
  ND2M1S U132 ( .A(n38), .B(n17), .Z(n20) );
  OAI21M1S U133 ( .A1(n17), .A2(n38), .B(n20), .Z(n18) );
  MAOI22M1SA U134 ( .A1(n19), .A2(n18), .B1(n19), .B2(n18), .Z(N201) );
  MAOI222M1SA U135 ( .A(add_regs[72]), .B(n126), .C(n20), .Z(n37) );
  NR2M2S U136 ( .A(add_regs[70]), .B(n37), .Z(n133) );
  MAOI22M1SA U137 ( .A1(add_regs[71]), .A2(n133), .B1(add_regs[71]), .B2(n133), 
        .Z(N203) );
  INVM1S U138 ( .A(add_regs[79]), .Z(n150) );
  ND2M1S U139 ( .A(add_regs[75]), .B(n150), .Z(n149) );
  ND2M1S U140 ( .A(intadd_2_n1), .B(n149), .Z(n22) );
  OAI21M1S U141 ( .A1(intadd_2_n1), .A2(n149), .B(n22), .Z(n21) );
  MAOI22M1SA U142 ( .A1(add_regs[76]), .A2(n21), .B1(add_regs[76]), .B2(n21), 
        .Z(N217) );
  NR2M1S U143 ( .A(add_regs[76]), .B(n22), .Z(n158) );
  INVM1S U144 ( .A(add_regs[77]), .Z(n157) );
  ND2M1S U145 ( .A(n158), .B(n157), .Z(n156) );
  NR2M1S U146 ( .A(add_regs[78]), .B(n156), .Z(n40) );
  MAOI22M1SA U147 ( .A1(add_regs[79]), .A2(n40), .B1(add_regs[79]), .B2(n40), 
        .Z(N220) );
  AN2M1S U148 ( .A(order[70]), .B(order[43]), .Z(intadd_35_B_1_) );
  AN2M1S U149 ( .A(order[74]), .B(order[106]), .Z(intadd_22_B_1_) );
  AN2M1S U150 ( .A(order[113]), .B(order[137]), .Z(intadd_27_B_1_) );
  AN2M1S U151 ( .A(order[130]), .B(order[139]), .Z(n136) );
  AN2M1S U152 ( .A(n135), .B(n134), .Z(intadd_0_A_17_) );
  AN2M1S U153 ( .A(shift_regs[160]), .B(shift_regs[8]), .Z(intadd_14_CI) );
  AN2M1S U154 ( .A(shift_regs[152]), .B(shift_regs[16]), .Z(intadd_13_CI) );
  AN2M1S U155 ( .A(shift_regs[144]), .B(shift_regs[24]), .Z(intadd_12_CI) );
  AN2M1S U156 ( .A(shift_regs[136]), .B(shift_regs[32]), .Z(intadd_11_CI) );
  AN2M1S U157 ( .A(shift_regs[128]), .B(shift_regs[40]), .Z(intadd_10_CI) );
  AN2M1S U158 ( .A(shift_regs[168]), .B(shift_regs[0]), .Z(intadd_15_CI) );
  AN2M1S U159 ( .A(shift_regs[120]), .B(shift_regs[48]), .Z(intadd_9_CI) );
  AN2M1S U160 ( .A(shift_regs[112]), .B(shift_regs[56]), .Z(intadd_8_CI) );
  AN2M1S U161 ( .A(shift_regs[104]), .B(shift_regs[64]), .Z(intadd_7_CI) );
  AN2M1S U162 ( .A(shift_regs[96]), .B(shift_regs[72]), .Z(intadd_6_CI) );
  AN2M1S U163 ( .A(shift_regs[88]), .B(shift_regs[80]), .Z(intadd_5_CI) );
  AN2M1S U164 ( .A(add_regs[9]), .B(N101), .Z(intadd_16_CI) );
  AO21M1SA U165 ( .A1(add_regs[30]), .A2(n23), .B(n24), .Z(N124) );
  INVM1S U166 ( .A(n24), .Z(n25) );
  OA21M1SA U167 ( .A1(add_regs[31]), .A2(n25), .B(add_regs[32]), .Z(N126) );
  AO21M1SA U168 ( .A1(N127), .A2(n89), .B(n26), .Z(N128) );
  AO21M1SA U169 ( .A1(add_regs[36]), .A2(n82), .B(n81), .Z(n27) );
  MAOI22M1SA U170 ( .A1(add_regs[37]), .A2(n28), .B1(add_regs[37]), .B2(n28), 
        .Z(n29) );
  INVM1S U171 ( .A(N127), .Z(n92) );
  INVM1S U172 ( .A(add_regs[34]), .Z(n91) );
  NR2M1S U173 ( .A(n92), .B(n91), .Z(n90) );
  NR2M1S U174 ( .A(add_regs[37]), .B(add_regs[39]), .Z(n74) );
  ND2M1S U175 ( .A(add_regs[37]), .B(add_regs[39]), .Z(n73) );
  ND2B1M1S U176 ( .NA(n74), .B(n73), .Z(n71) );
  MAOI22M1SA U177 ( .A1(n71), .A2(n88), .B1(n71), .B2(n88), .Z(n31) );
  OA21M1SA U178 ( .A1(n146), .A2(intadd_30_B_1_), .B(n145), .Z(N146) );
  AO21M1SA U179 ( .A1(add_regs[46]), .A2(n147), .B(n32), .Z(N154) );
  INVM1S U180 ( .A(n32), .Z(n33) );
  OA21M1SA U181 ( .A1(add_regs[47]), .A2(n33), .B(add_regs[48]), .Z(N156) );
  OA21M1SA U182 ( .A1(intadd_32_B_0_), .A2(intadd_32_A_1_), .B(n34), .Z(N159)
         );
  INVM1S U183 ( .A(add_regs[51]), .Z(n98) );
  OAI21M1S U184 ( .A1(add_regs[49]), .A2(add_regs[50]), .B(intadd_32_A_1_), 
        .Z(n35) );
  ND2M1S U185 ( .A(n98), .B(n35), .Z(intadd_32_CI) );
  MAOI222M1SA U186 ( .A(n104), .B(n102), .C(n101), .Z(n36) );
  ND2M1S U187 ( .A(add_regs[55]), .B(n36), .Z(n103) );
  OA21M1SA U188 ( .A1(add_regs[55]), .A2(n36), .B(n103), .Z(N170) );
  OA21M1SA U189 ( .A1(n120), .A2(n114), .B(n119), .Z(N175) );
  OA21M1SA U190 ( .A1(n131), .A2(n125), .B(n130), .Z(N191) );
  AO21M1SA U191 ( .A1(n37), .A2(add_regs[70]), .B(n133), .Z(N202) );
  INVM1S U192 ( .A(N189), .Z(n128) );
  INVM1S U193 ( .A(add_regs[65]), .Z(n127) );
  OA21M1SA U194 ( .A1(add_regs[71]), .A2(n39), .B(n38), .Z(intadd_3_A_6_) );
  INVM1S U195 ( .A(N206), .Z(intadd_2_A_3_) );
  NR2M1S U196 ( .A(add_regs[73]), .B(intadd_2_A_3_), .Z(intadd_2_CI) );
  AO21M1SA U197 ( .A1(add_regs[73]), .A2(intadd_2_A_3_), .B(intadd_2_CI), .Z(
        N208) );
  AO21M1SA U198 ( .A1(add_regs[78]), .A2(n156), .B(n40), .Z(N219) );
  INVM1S U199 ( .A(add_regs[75]), .Z(intadd_2_B_1_) );
  INVM1S U200 ( .A(add_regs[76]), .Z(intadd_2_B_2_) );
  AOI21B20M1S U201 ( .NA1(order[70]), .NA2(order[43]), .B(intadd_35_B_1_), .Z(
        n43) );
  AOI21B20M1S U202 ( .NA1(order[74]), .NA2(order[106]), .B(intadd_22_B_1_), 
        .Z(n48) );
  AN2M1S U203 ( .A(order[108]), .B(order[132]), .Z(n139) );
  AN2M1S U204 ( .A(order[111]), .B(order[135]), .Z(n138) );
  AN2M1S U205 ( .A(order[112]), .B(order[136]), .Z(n137) );
  AN2M1S U206 ( .A(order[129]), .B(order[138]), .Z(n69) );
  AOI21B20M1S U207 ( .NA1(order[129]), .NA2(order[138]), .B(n69), .Z(n64) );
  ND2M1S U208 ( .A(intadd_16_n1), .B(add_regs[14]), .Z(n141) );
  OA21M1SA U209 ( .A1(intadd_16_n1), .A2(add_regs[14]), .B(n141), .Z(N110) );
  OA21M1SA U210 ( .A1(intadd_25_A_0_), .A2(n70), .B(n143), .Z(N116) );
  AOI21B20M1S U211 ( .NA1(shift_regs[168]), .NA2(shift_regs[0]), .B(
        intadd_15_CI), .Z(N1) );
  AOI21B20M1S U212 ( .NA1(shift_regs[160]), .NA2(shift_regs[8]), .B(
        intadd_14_CI), .Z(N10) );
  AOI21B20M1S U213 ( .NA1(shift_regs[152]), .NA2(shift_regs[16]), .B(
        intadd_13_CI), .Z(N19) );
  AOI21B20M1S U214 ( .NA1(shift_regs[144]), .NA2(shift_regs[24]), .B(
        intadd_12_CI), .Z(N28) );
  AOI21B20M1S U215 ( .NA1(shift_regs[136]), .NA2(shift_regs[32]), .B(
        intadd_11_CI), .Z(N37) );
  AOI21B20M1S U216 ( .NA1(shift_regs[128]), .NA2(shift_regs[40]), .B(
        intadd_10_CI), .Z(N46) );
  AOI21B20M1S U217 ( .NA1(shift_regs[120]), .NA2(shift_regs[48]), .B(
        intadd_9_CI), .Z(N55) );
  AOI21B20M1S U218 ( .NA1(shift_regs[112]), .NA2(shift_regs[56]), .B(
        intadd_8_CI), .Z(N64) );
  AOI21B20M1S U219 ( .NA1(shift_regs[104]), .NA2(shift_regs[64]), .B(
        intadd_7_CI), .Z(N73) );
  AOI21B20M1S U220 ( .NA1(shift_regs[96]), .NA2(shift_regs[72]), .B(
        intadd_6_CI), .Z(N82) );
  AOI21B20M1S U221 ( .NA1(shift_regs[88]), .NA2(shift_regs[80]), .B(
        intadd_5_CI), .Z(N91) );
  INVM1S U222 ( .A(add_regs[40]), .Z(n94) );
  INVM1S U223 ( .A(add_regs[38]), .Z(n78) );
  NR2M1S U224 ( .A(n94), .B(n78), .Z(intadd_1_B_9_) );
  AOI21M1S U225 ( .A1(n94), .A2(n78), .B(intadd_1_B_9_), .Z(intadd_1_A_8_) );
  ND2M1S U226 ( .A(add_regs[40]), .B(add_regs[36]), .Z(n72) );
  OAI21M1S U227 ( .A1(n74), .A2(n72), .B(n73), .Z(intadd_1_B_8_) );
  OAI21M1S U228 ( .A1(add_regs[40]), .A2(add_regs[36]), .B(n72), .Z(n77) );
  OA21M1SA U229 ( .A1(n74), .A2(n88), .B(n73), .Z(n76) );
  INVM1S U230 ( .A(n75), .Z(intadd_1_B_7_) );
  INVM1S U231 ( .A(n79), .Z(intadd_1_A_6_) );
  INVM1S U232 ( .A(add_regs[39]), .Z(n86) );
  INVM1S U233 ( .A(n80), .Z(n85) );
  AOI21M1S U234 ( .A1(n82), .A2(add_regs[37]), .B(n81), .Z(n84) );
  INVM1S U235 ( .A(n83), .Z(intadd_1_B_5_) );
  INVM1S U236 ( .A(n87), .Z(intadd_1_A_4_) );
  NR2M1S U237 ( .A(n88), .B(n91), .Z(intadd_1_B_1_) );
  AOI21M1S U238 ( .A1(n88), .A2(n91), .B(intadd_1_B_1_), .Z(intadd_1_B_0_) );
  AOI21M1S U239 ( .A1(n92), .A2(n91), .B(n89), .Z(intadd_1_CI) );
  AOI21M1S U240 ( .A1(n92), .A2(n91), .B(n90), .Z(intadd_1_B_2_) );
  INVM1S U241 ( .A(intadd_1_n1), .Z(n93) );
  NR2M1S U242 ( .A(n94), .B(n93), .Z(N141) );
  AOI21M1S U243 ( .A1(n94), .A2(n93), .B(N141), .Z(N140) );
  OAI21M1S U244 ( .A1(n100), .A2(intadd_31_CI), .B(n95), .Z(intadd_31_A_3_) );
  INVM1S U245 ( .A(add_regs[52]), .Z(n96) );
  ND2M1S U246 ( .A(n101), .B(n96), .Z(intadd_31_B_3_) );
  OAI21M1S U247 ( .A1(n96), .A2(n101), .B(intadd_31_B_3_), .Z(intadd_31_A_2_)
         );
  INVM1S U248 ( .A(n97), .Z(intadd_31_B_2_) );
  INVM1S U249 ( .A(n99), .Z(intadd_31_A_1_) );
  INVM1S U250 ( .A(intadd_31_SUM_0_), .Z(intadd_32_A_3_) );
  ND2M1S U251 ( .A(add_regs[50]), .B(n100), .Z(intadd_32_B_2_) );
  OAI21M1S U252 ( .A1(add_regs[50]), .A2(n100), .B(intadd_32_B_2_), .Z(
        intadd_32_B_1_) );
  INVM1S U253 ( .A(intadd_32_n1), .Z(intadd_31_B_1_) );
  AOI211M1S U254 ( .A1(n102), .A2(n101), .B(n104), .C(intadd_31_CI), .Z(N172)
         );
  AOI21M1S U255 ( .A1(n104), .A2(n103), .B(N172), .Z(N171) );
  INVM1S U256 ( .A(intadd_32_SUM_3_), .Z(N165) );
  INVM1S U257 ( .A(intadd_32_SUM_2_), .Z(N164) );
  INVM1S U258 ( .A(intadd_32_SUM_1_), .Z(N163) );
  INVM1S U259 ( .A(intadd_32_SUM_0_), .Z(N162) );
  OAI21M1S U260 ( .A1(n123), .A2(n106), .B(n105), .Z(intadd_4_A_6_) );
  INVM1S U261 ( .A(add_regs[61]), .Z(n107) );
  ND2M1S U262 ( .A(n107), .B(n106), .Z(intadd_4_B_6_) );
  OAI21M1S U263 ( .A1(n106), .A2(n107), .B(intadd_4_B_6_), .Z(intadd_4_A_5_)
         );
  ND2M1S U264 ( .A(n107), .B(n108), .Z(intadd_4_B_5_) );
  OAI21M1S U265 ( .A1(n108), .A2(n107), .B(intadd_4_B_5_), .Z(intadd_4_A_4_)
         );
  INVM1S U266 ( .A(add_regs[59]), .Z(n110) );
  ND2M1S U267 ( .A(n110), .B(n108), .Z(intadd_4_B_4_) );
  OAI21M1S U268 ( .A1(n108), .A2(n110), .B(intadd_4_B_4_), .Z(intadd_4_A_3_)
         );
  INVM1S U269 ( .A(n109), .Z(intadd_4_B_3_) );
  INVM1S U270 ( .A(n111), .Z(intadd_4_A_2_) );
  INVM1S U271 ( .A(add_regs[57]), .Z(n115) );
  INVM1S U272 ( .A(n112), .Z(intadd_4_B_2_) );
  INVM1S U273 ( .A(n113), .Z(intadd_4_A_1_) );
  NR2M1S U274 ( .A(add_regs[62]), .B(n115), .Z(intadd_4_B_1_) );
  AOI21M1S U275 ( .A1(add_regs[62]), .A2(n115), .B(intadd_4_B_1_), .Z(
        intadd_4_B_0_) );
  INVM1S U276 ( .A(intadd_4_B_4_), .Z(n116) );
  AOI31M1S U277 ( .A1(n116), .A2(n115), .A3(n114), .B(N173), .Z(n117) );
  NR2M1S U278 ( .A(add_regs[61]), .B(n117), .Z(intadd_4_CI) );
  AOI21M1S U279 ( .A1(n117), .A2(add_regs[61]), .B(intadd_4_CI), .Z(N178) );
  AOI21M1S U280 ( .A1(add_regs[59]), .A2(n119), .B(n118), .Z(N176) );
  AOI21M1S U281 ( .A1(add_regs[57]), .A2(N173), .B(n120), .Z(N174) );
  AOI21M1S U282 ( .A1(n123), .A2(n122), .B(n121), .Z(N188) );
  INVM1S U283 ( .A(add_regs[70]), .Z(n124) );
  NR2M1S U284 ( .A(add_regs[67]), .B(n124), .Z(intadd_3_B_6_) );
  AOI21M1S U285 ( .A1(add_regs[67]), .A2(n124), .B(intadd_3_B_6_), .Z(
        intadd_3_A_5_) );
  NR2M1S U286 ( .A(add_regs[66]), .B(n126), .Z(intadd_3_B_5_) );
  AOI21M1S U287 ( .A1(add_regs[66]), .A2(n126), .B(intadd_3_B_5_), .Z(
        intadd_3_A_4_) );
  ND2M1S U288 ( .A(n124), .B(n125), .Z(intadd_3_A_2_) );
  OAI21M1S U289 ( .A1(n125), .A2(n124), .B(intadd_3_A_2_), .Z(intadd_3_A_1_)
         );
  ND2M1S U290 ( .A(n126), .B(n127), .Z(intadd_3_B_1_) );
  OAI21M1S U291 ( .A1(n127), .A2(n126), .B(intadd_3_B_1_), .Z(intadd_3_B_0_)
         );
  OAI21M1S U292 ( .A1(add_regs[68]), .A2(n129), .B(n128), .Z(intadd_3_CI) );
  INVM1S U293 ( .A(intadd_3_SUM_6_), .Z(N200) );
  INVM1S U294 ( .A(intadd_3_SUM_5_), .Z(N199) );
  INVM1S U295 ( .A(intadd_3_SUM_4_), .Z(N198) );
  INVM1S U296 ( .A(intadd_3_SUM_3_), .Z(N197) );
  INVM1S U297 ( .A(intadd_3_SUM_2_), .Z(N196) );
  INVM1S U298 ( .A(intadd_3_SUM_1_), .Z(N195) );
  INVM1S U299 ( .A(intadd_3_SUM_0_), .Z(N194) );
  AOI21M1S U300 ( .A1(add_regs[67]), .A2(n130), .B(n129), .Z(N192) );
  AOI21M1S U301 ( .A1(add_regs[65]), .A2(N189), .B(n131), .Z(N190) );
  AOI21B10M1S U302 ( .NA2(add_regs[71]), .A1(n133), .B(n132), .Z(N204) );
  AOI21B20M1S U303 ( .NA1(n135), .NA2(n134), .B(intadd_0_A_17_), .Z(
        intadd_26_A_3_) );
  AOI21B20M1S U304 ( .NA1(order[130]), .NA2(order[139]), .B(n136), .Z(
        intadd_26_A_1_) );
  AOI21B20M1S U305 ( .NA1(order[113]), .NA2(order[137]), .B(intadd_27_B_1_), 
        .Z(intadd_34_A_1_) );
  AOI21B20M1S U306 ( .NA1(order[112]), .NA2(order[136]), .B(n137), .Z(
        intadd_17_A_1_) );
  AOI21B20M1S U307 ( .NA1(order[111]), .NA2(order[135]), .B(n138), .Z(
        intadd_18_A_1_) );
  AOI21B20M1S U308 ( .NA1(order[108]), .NA2(order[132]), .B(n139), .Z(
        intadd_21_A_1_) );
  INVM1S U309 ( .A(add_regs[15]), .Z(n140) );
  NR2M1S U310 ( .A(n141), .B(n140), .Z(N112) );
  AOI21M1S U311 ( .A1(n141), .A2(n140), .B(N112), .Z(N111) );
  AOI21B20M1S U312 ( .NA1(add_regs[9]), .NA2(N101), .B(intadd_16_CI), .Z(N103)
         );
  INVM1S U313 ( .A(add_regs[29]), .Z(intadd_25_B_4_) );
  INVM1S U314 ( .A(add_regs[28]), .Z(intadd_25_B_3_) );
  INVM1S U315 ( .A(add_regs[26]), .Z(intadd_25_A_1_) );
  OAI21M1S U316 ( .A1(N115), .A2(n142), .B(intadd_25_B_2_), .Z(intadd_25_CI)
         );
  INVM1S U317 ( .A(intadd_25_SUM_4_), .Z(N123) );
  INVM1S U318 ( .A(intadd_25_SUM_3_), .Z(N122) );
  INVM1S U319 ( .A(intadd_25_SUM_2_), .Z(N121) );
  INVM1S U320 ( .A(intadd_25_SUM_1_), .Z(N120) );
  INVM1S U321 ( .A(intadd_25_SUM_0_), .Z(N119) );
  AOI21M1S U322 ( .A1(add_regs[26]), .A2(n143), .B(n142), .Z(N117) );
  INVM1S U323 ( .A(add_regs[43]), .Z(intadd_30_B_2_) );
  INVM1S U324 ( .A(add_regs[41]), .Z(intadd_30_B_0_) );
  OAI21M1S U325 ( .A1(N144), .A2(n144), .B(intadd_30_B_3_), .Z(intadd_30_CI)
         );
  INVM1S U326 ( .A(intadd_30_SUM_3_), .Z(N152) );
  INVM1S U327 ( .A(intadd_30_SUM_2_), .Z(N151) );
  INVM1S U328 ( .A(intadd_30_SUM_1_), .Z(N150) );
  INVM1S U329 ( .A(intadd_30_SUM_0_), .Z(N149) );
  AOI21M1S U330 ( .A1(add_regs[43]), .A2(n145), .B(n144), .Z(N147) );
  AOI21M1S U331 ( .A1(add_regs[41]), .A2(N144), .B(n146), .Z(N145) );
  OAI21M1S U332 ( .A1(intadd_30_n1), .A2(n148), .B(n147), .Z(N153) );
  OAI21M1S U333 ( .A1(add_regs[75]), .A2(n150), .B(n149), .Z(intadd_2_A_7_) );
  INVM1S U334 ( .A(add_regs[78]), .Z(n151) );
  ND2M1S U335 ( .A(add_regs[74]), .B(n151), .Z(intadd_2_B_7_) );
  OAI21M1S U336 ( .A1(add_regs[74]), .A2(n151), .B(intadd_2_B_7_), .Z(
        intadd_2_A_6_) );
  INVM1S U337 ( .A(n152), .Z(intadd_2_B_6_) );
  INVM1S U338 ( .A(n153), .Z(intadd_2_A_5_) );
  INVM1S U339 ( .A(n154), .Z(intadd_2_B_5_) );
  INVM1S U340 ( .A(n155), .Z(intadd_2_A_4_) );
  ND2M1S U341 ( .A(add_regs[77]), .B(intadd_2_B_1_), .Z(intadd_2_B_4_) );
  INVM1S U342 ( .A(add_regs[74]), .Z(intadd_2_B_0_) );
  OAI21M1S U343 ( .A1(add_regs[77]), .A2(intadd_2_B_1_), .B(intadd_2_B_4_), 
        .Z(intadd_2_B_3_) );
  OAI21M1S U344 ( .A1(n158), .A2(n157), .B(n156), .Z(N218) );
  INVM1S U345 ( .A(intadd_2_SUM_7_), .Z(N216) );
  INVM1S U346 ( .A(intadd_2_SUM_6_), .Z(N215) );
  INVM1S U347 ( .A(intadd_2_SUM_5_), .Z(N214) );
  INVM1S U348 ( .A(intadd_2_SUM_4_), .Z(N213) );
  INVM1S U349 ( .A(intadd_2_SUM_3_), .Z(N212) );
  INVM1S U350 ( .A(intadd_2_SUM_2_), .Z(N211) );
  INVM1S U351 ( .A(intadd_2_SUM_1_), .Z(N210) );
  INVM1S U352 ( .A(intadd_2_SUM_0_), .Z(N209) );
endmodule
